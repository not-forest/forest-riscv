`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MX91U1xqdDZcPCpmcsBSmjipgmG1OTfore0cfYMDQr3pZ6ENndD53F996zXgdori
2W3jy4q9Mm+TqH+CdktNFEEYMpLcIUeuBEQudkvpQBqSmQ/3GuH63FszgSBlODjS
qHTL3m1gkwu/ebQ8jiXwPa5J8ftXgjSuD69oHeb50b8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21696)
fzMX5mfNZcFPOO1Nq5AkZBrSMBVk57NVqFFAUfoOk8Usm3pQLiealJd+fecUODel
C9FbYVJWIphgrnzwL5F2cEmxJxUFcf6PACErKypj5oeE05OtHTcVvgMTbQu5/rnx
zmW5H4HImfrqQlpd2Uvy832tSxNIekRrtQTp4l10Tk6Y9LphuTnypZzZU8R/vTrI
JieZllihXphgqSELonkyWl/YYBjXGcdIQGw0t2VhaBWPLs3J1twYOL3w7VkJyZnt
jbnK46WwRqkGOndAGm8EOPhYEFt+lvTicDn116oyHYPyFWfEaUAdIvTk/0rZ+U/X
rf8dGhs6DEhpju2y3a35g36MEUPT2mjoSx6rWnnwOp23zpXTU8H4bJ0hCuqyv9Np
dHHpFFAmaHpxjq5pxwGqNqniSC9y4JH03/JIfZSIBL6o7OTl4h7E0Pk6TIx4cb+w
ov7J57bp4I1TyCI6oVZzJpNodGSecHdjDj0K3vPSTDcpX1Q6JwGcu8NvbGQ26spO
gbSX2lp1gEmhJWTRULCThghi55IaNvvRs/U89yRDbxpLMPWbKsa1KQnX3dUi8pWM
t9JPJgWFBY1BQHgAp2HFsKaLpuhRXA4Kaciths3Gi9wUIyaaniSb0AUcA0ci9q+0
GiIh3V642XqsozBvCcMB25KuVf0WSaUeHf8ka1T4fo7cwdHGSjy3JPx7P4S9pYwU
tZOtE2t5FX8cXo58jAPrfOlL7eLqrJtdDxSeXZPbwUfcE4KtInxKhY/WNeCF5gJw
3t+SQBTdYzyQzVuw41zZn+d1EYKcZlIediIRXJbM3mwp6E9uH6yqEbp9IsXq7rZh
hi88OYGAbc6Yn6F9OUB8quXXBzhKaVzzXn0wI+nwxUVeUuoa2QEC64UAh7BCZG+4
gnlATOxIxVhQ8k7tC743TS29+COckL8b7l+/UEC9QCIX17Jr0vGmno0guw9HyzhK
/0U5RgSaLRZaJb9BW/S1LeOapNAH7vDjr1iOeEih+GCXmkN5kjpgoFZpX+X/i0MB
aIQRYNUAXI0Q/My6MqNllTu5hvlrDeOmzhDrbW/W5ps0w5UIW+Qnt3gJ2PsU/CAq
hzdSavmXoieYXk5dUSC4MPqmb1JqhhF4+Z08ilvJRzQqu3wFUBNEFyrf8psA/b2z
hV4HvfYoT6UWjJr3334YxtaKCKfq6KBMHZac87hQ5/2LqqZwcLzkyyKEb7w899eg
mhpaqVcoOhCuFPMsmzhjjmAJCwL1948YJJ9Q7TfvRYpt4GSdVzSAT1S7rlyImhjx
WhegdIqjA6411A76Bqaw0zIp0yoIXA3yH4tguWQZbuWlP4DaTLzRCtK41mXfAnRy
KkceWhG46KoQ4/ieWiFJo6EbAqm+xcak4AwipqNWRP7wQLyJ39PlNaPz0/AegfH1
9KuUzEvqYj2iHgDDW9oFdqTw0HorU2TGhusYa2PtuT3BCMz01B88yiuKO7WtGBoH
D2m8WNmx2y3BJ8l8hJKUJcnReXKPRgHFPbsQwxUedTXVWMHVx6Z4ghKSrxRgZSiE
y/+B9eMoHBkVi/D42skxGO8Mq3QHzJnGaCRuyYm1/qflAU7i2rP2LtFywf23r/sO
JtRqEoBKr3FZ3nu1j7fY8hhr6Lommjc4lBGzdJBkgYwbOuedIaUOD4cRXWPLpJMT
GV9KwIPvOiSyNWQF75WZ2GRDt4MNbiCcY1x26VxnD/pPq09ggLvrUomP8r9JLWkt
p/wb0dMK5zeVDT78/w1x3ZNftWAC6WvmZy49a0OtCJVnukDJIBH4kAQagadPwdfj
qiIbktM1SrWzWvZubtUby5KoNZrjdoFP14k0LQaxBCSmx+mU2zHvwHmlAz0ECn9A
sXHx+aXCHGC5wxcuLI6LmyyIQbCvoHqPd4wFpMXcnBrVArQ+P7y1+ITwzfgK0Yco
r/jSe/KhaNf9lZfTPUQ830pCtWzKgC0DWUuo3kncHZRG7oESlGd+zTtMuqW9ICGh
kcXDZKM2OAJwSsLeqtVh0Od9QuaQxCSuJyDTS1yccq9cncudrPXYlKUFYZ69tieH
0vM0UyqAt9L7gH8T/AxwAVWcF+dLhI5d6VVNvo+MJLEd0vzzgl4YfVS+dqqc3EqG
4uuu+YaXeS+lt+oV7P9WEiK9YZXVxvKF2Ck7sb+g81KQ5vLQy1o2FgaktsZDuFMG
WPCo08kRail9p/ZHGdMPegOIaY0Pi+HA6Q+o1Ouax2A5ONXmG///SeyBSTXYPSJO
2TQGhiYhG4YELQVjDt1nKin/x1VxthJLNk/o87DEzCccl9Np1AhLrnEM200AHIS3
G1Em5nkMoQd7/OA8VeKNgMLqwysEleHvX/2XDtEX+JV3Jk5gzNFeyGY5bwcH1y+l
4r0fICwnBSrnBWUpaqD8PbqZERC06sohuGM03GIrtQpVDrQyhkSArXEA4HC5OFI0
UKwZzPA23m/L2wIrVEug5KVsXgJFtDYzv4+fR0dqRI9gBfOQAh3i7rW/zqnMeR0/
QWoAnKnATE03hxl8hsDpJ3IzFr/sB8lOFMTcj60qcXi3Zjibh0OgmHv1in7OCOL+
DJfGFgnmizcgmuArRl3INBPeRxqW1X0jAmaB2jWlc2IFU+CTE9kpkEbmzJGasxrL
IOvBHJgSh8HgV7vZsaSWXSQYgMA31zJLV6klAMMKQnFwoGeC1qgXUGdi4vyVe08h
O+vu7gT4p1H8x37JRF8Nl70rRpj87sTvEKB6CHvJr2A/IeY/yW0HFZeMT+7fDRKH
MykIIwXQPrq7sdXr95TI/cuNvJfLjdseuHzAmaM1AIR4EyH7Q8YbLZToU9bCPgpe
PBr7CipDiGKB+NEd6DeU19HkQ8zWHTEqiWDR6FrehmTaCkqZQvuokm80q6SCCigt
G0wuBsph7+MRDoRfnZ1FMyHIIJ2k44oeiEBg/VAXUIyUycbFiMMcNBdT4+ClQCNn
DKVOMgLV0wl7xu3OmDu5Jpj3xLaQDlMXIpufEY8TGSjuhUB1AuLGYLVo4rraLvyh
LYU5IMnzbQxGsFfXkpvpleZKwFLF0OEbbvHcRTTW5CQPhQHhZ9RlxU57+HWxpuWU
63uZXbx79MAnhnZ06XqD187A6ZYEXPK/ToBWgq6NfDcA5zZJD+5Di427jCgPq/eR
ATpDJlfWNmw/XGSzuMh6fDIdlUsIjUxGhDo8EFQEmRACFYvkHQcsJoztr5+7UjRG
Zk6L+mDoBn5cPg0D6I/54fRdwDJoydHwoY8NIY0oxDonJ4nPMeHYH9HMwlD0vCIu
RXNZGwVLQZ4g0tQUJk2lD+7Dz/NzUfJHniqC5Nd6eHIfPy/Z5I1O20M2FCXfyh/L
vxYy9P4P3xxOLi2piOwS3ETGvGVmTwxcnfQglvk2Y0reCHG2h/xFO9XYcBAGc3+w
um3chE/QAoCnsy72Jssgvyx1E5J/n3WnL+BYCBcznO3aToxRfhV8+xcCZgmkGUpk
gmWhBhrHgtwslJxqvqn6KY667ZVU2LTfFLgb1AbirWPrvXDczRAYbGWEoLOYH0RH
OofoUgurGPyobKBvyrqkOSHUk08lGWtjPPnVRsMXh7iyrvt320A7SPavcCEb6rJL
XalaazGAqBOKPPg1sYEFHoZ9Go+d0FC5saZDzTE5wcr9bi9Ix7onLEpffEfDkDnE
YOAlpbmPgBF9Z0gL10pyM/HcPBpfCiE6IJ1Wzm/k22pwELBRBxcDuHfKLZ8sdP6+
fiBovqqV32ZATImsWVuiuPZfOJ9CrdATKJnfT5lD9ruOc5ZXJp9DsUCnJRow/ZLI
did30Calp5zH4FN52l8qYa6HLsC0A5HtRSF9OczCrPjfYWi+DQUog/KtDSDUpPkJ
K1fe82O8Qq/eoBENdcW/QDbcZUu+UUp5S8Tzsng85VyWXkW7fLXJQSuFN62wisNi
YDxo7D6rpzmDshZ+uOPcgEDx5M5PXTWkp+VH9ZELzteyeGwU/uA2kF/fyrU3A8HB
LiYAAbi34Fe17WcT/Nsn39KjUGmr/sn5RwTeYvYLExfHxZ7TEKYDZbdrL4q671R4
VjxJqqot26JIHsZGYV8CkBQopWkmLHMt7PeiTIVtD2+WzGJWABq0OYAfB3rIvYyo
ODXHxU9u+ZWuXq12dHz9mmfxmlEMNJCYYT5cOte4z+dGAN3iOu9Ez8GnUYBP4sUa
jyGeQvVkLpC2oeXKo0FyeV5XO17IiQRXGoDCdwx9dW5KEEodNwjzraf0w1t8wZSB
0u9kqsOU4Ci+2JZEU9Cb09H1NFmLILgL4p0BGLN2L9JvfR2VVBEuGJqwli7ZKOar
3cLM5TmQHfPYEkLSMX5OJWtv2Iih2Y7ono/ldPNaS4UltvqjbPnUvO8E3kVg+ePl
p1PlY9qciit+2DRr/97tjYUpsi8sO8BvOvddJpSvQdd7cuBaAo2UvJuZYuOS+e8u
IvF35vzvgVGzWkso/y23ef5iTNBmQIwdU2lzD5DXvHU7rYBVcaqGqoj7ZflapXJv
Ivq5qbo274nENxYUFQWrtxPuf+qTYd77SROCzMPP7xbUVAk1ATy3tl85sjsLNgk6
7b2u/17p+iySIgcatI3x6vIkOlRcyiiLuFm3vVtOFdHScSHExvJVUt2Uk7VUQ6FK
0Czet0ihkgcswheSVa9vQf1C9aeloOQFlM0Lk3ZEWjPxaBkHyzL8KS2VCGj5QGkD
orWMFx8FAuOqjKkpBqY5WMl6Edln7hakcri/CAj8LwP2WBNH/901XDghmd2sTkYb
sucEY+tbYZ999NpPeZGEV+iHFp6nv7P+9r2z6mnyI6g62XFHN3UvlAGKQ89KVYHS
qo/8uHcjS5raOr3fy6sS9/AkbW/fllGUuPIyurNsjgJGWSnBlossCDWDIrJ9KhRC
iJ7VQtIUl9Ew4hjavqpCWZPhutcP1IZf0pf8ufSTxGgfGF362mbFAdQ8Sl0U6PNn
p5ntYjVnW4X+jwtMzQiQMZ2vbpeOjfiE92pBQ3lLR6+IpXJS0aLdgZRxB+C62YQr
molouTK8QkOr/gPpxTIKidZGwKLD6lY/NMO1WOOvoKYQxToWeZ9KdPwypSUUxHZ4
x/0cSSB3CrSoy/34aUlrxhMZiXLojIO6xy8szEO6bfhmEkGJh40AhRkr3CROwMTH
ZvQSMV3wA14lmTpPci6/ByXDJZ+mbZNkazt2QCE31hSFKrLjjQC1EdRni3vA4SBy
gcSOoHowg0YlyaSLFdW1I1uUzsCisYu2XmQjq4UqTLV5MVzh4/elXP+JO5j8gWul
pMzPfKTFCdLZe2Ew4CAqNGSpRLI7X6PykpA1w0OF+DzP0qd/koiiXn2nJUH+JcRh
owSIlauZdGd0AkTseBj2D81pPHEUtTRCO8h7FmbLjWC3YMx5Es2HdNdrJowSgFn7
7QRYj7oF+dsHlXkc8U/2/asuGSiHhMDMk6UpGy9efdjP/+8ouVkq1SA4WXZTFLZg
Iijelb5EY+NwOPniU8RC63tCQtmy9/ZE/YG7LPDqu3TnmdEU9WL6K4RYIK8nbgW4
babLGKjm4Oyi3yMR2WjJNmCK8bqochvmt4KqVHt4hHlILyENhbyl//5Mq3dluROU
EUkiq7OPWXf+EPN8eevUPMbpxsXNNrYJ5leGSvrrNvEiTlRQOnNTqvblq1QLTfxF
NthGd0KJFEEXAbLpdZjkLIGya0y1qWlyH31HAoMrIOCz8GMn/IfEQ9ved6YIzpf1
nOtFC+OhUnMLX/3V+rliPp3YhNAhz+xxA3VwVm2oRFH0oyyS/ET+IDqagy3m8bJd
KorNn5f5katra2IG9yeqXf1UbGg9v28EJeEB2JSjop/KeRrzhI2mlU3i0OWbaNm6
2W9t6XVUwSAon8aBT8HS9I5WDNzhScGbI0HWZ1lYdLkX4pJ3RAtRiBctSQr2hUvk
GOJF1WwAHGJVWFNUqUtDk1MfgsWBCDem8Amimhh9f3kBqfl4yA/ubotSiPR6/9gk
mBzCJK2ZnBCpyrh6oGE7jugUyCV9WrDPnHw+Jc55BX0cDEPO7Q03sDOmSVqyi2R5
GR77kmw1ZPD29XTcGrieKhppMUuAx9o6VjYv/mjJoVYb9juOd9Xj/tJNtSdPFmIE
CKEmuz+AbljetKd66MJpfb9/3HbBHvmNmcx9AJ1eCz9wDJUHdzZt1TuulmJJTzf0
6J80JdcsgXUUs/wFJ6h8QVqTjnJPcoOdPfINMCqav28mTfAIlocPkwcxOKjIqEzq
Wxi7sv3SaB4BAil3LRtNlej5IU9nizdbVd55yswa2GR091TrH9/sv7K6pfpKKWKq
zMW8n5jh5f8C0KNSeil9zVXeKs/2+xGk/dFfF6Xkq/PFXQXW41CpmK9MoyHknGyE
g8BSqdAX6UZz7PnHP6mN6TM9lbmt4ureBqUrdAkFhIgUVVFlhBGVHZ69tOx+3lCU
G/WTSwhREq39/iy/TyN6zZexngw53FD7g3FxmWnqpobwIpgNbmIqREMWGs5M2gBP
2+hxoKQHwPfa8e3wJowd2LT4oDZCh1i0qY7qFfzSWDutEI0jI3GGq/sP75DY5RZY
bFzu7Ot4cGs4qRb2R+l58RivRDlW8bjXe0nuUJgjKg6+5tfa+TWStQaTWpd/oqwn
pUTJ2caecR+SpatKLlrO/2vkJWIeVkImMT4Jk+QgYHAxyzD25ZJX4rhC/Z5R3owd
SLLiBCkqW/Rjs7U6UPo1OvPyeH5rqlfcxtVWBjCMqJ3rhi4uREwv8VATx5hHRfN/
enOlv4GQYXpamAJKcLYf3X7oIYk7fewiWWHKS6XPFTC0HLdsm/mCSX2twQaJ8oCA
kcC+nGUFl/1WcJ2cCpw71R1UZeNOoW3tokDD7u9qzCSGxVQSL7PIzJgCHwo0gXyR
8UdZB3Bi7JhoMp4Lj/01ztk4vLE0jFy4+QJriJeTQtEFpHTKrKNmOrb5V2MTCLnU
+kRdroqjA8bWKbPZ5IhhB+gv1v8DqeylvOIcj825LN4A5GQTObSPXt6D1rzq4VJl
1SqRXKHYC4ADuFw0PBMwCMayMOpNwIvCNf+7abVccF+0W9um0SZ6W2aeqc4yYBgl
kFM6Oh59IQaMI6tJYmPYofNpjerENK2XLzDnbk1jfr5PtMLRO8kryxPuArCBsivv
eeT85yKJHm46/u4U/996DXSq78q2J/+r6vCJPg8mYhicVhy/hXKkXq5QjV6NFd6e
cthXHHdcQSK0sUvmDyJ4028uddwvEN1OY57JQCEQSn/7qutcSXrgd+4vxNWgTDFG
N0Q1N5LljW0Pa70vONe7ZYBjEqY/KLCfG/G21e5XQF3fssBk/er1g1Hq7sqq4NeB
SRju2P6Tr3l5pq8KOcKsh90m/uySbYJK0HkB7B3QRq90jN7mtzrnQnLZJ8ybK5uZ
Il/psPUYWqkhswaa0lujkw4pegSeHZOV+OmLttmWj+XdMS9b5yyYPmwfZWjdMbL5
k9DCNfkmMAf2Z+1Oy9qplo8bb+NfpQDfGhmdTEF+on7z/Ecw08D7IAaYVTcbCwvc
NBR7yCsJsuudBGQq4WG2/M2w8pp8kiVn5Rf9gZuWinjVl0iYGUTLdSgE++/5r+Q5
nToKbOcN8cTdw1rKy7hMiy0xv2MBKW4nQXaJhTWHWzBvOTp/S+AwCq8CM8S2POpf
z8jkfPc7bODlIkYBIFgNrDE1KSMBLG9tRBX6dD+jXeNdiZBouhG6tpqhVIIOd0+o
srBaSCyyF4WTdYdbVoZjWh0hlDr+yXLiA8jRjFgI3np+/p+CifkmmE0KSLlYDxvg
xRAe/qIGKJC4H/xDEwQX/laDEXRra7tf05eKag1NDZDJwwGq7BuvW0YA8B/y87D/
atmi55WfSNZXGfHA5oS8APDT4KCHjkltaAAVeLGmypMEgfRY4aMWqZQciGtuowni
6t61VPbP3uSZLy9lsAZd+4nAU+Vr3FxmQNoMlbDfHAcgKR6n3VJH5FDHiJ73K+uM
X92eFMpMXbNl6re3Ia55sXICZ+J3OG/vu5WDfrBxblwdMou2YBySHO+N0bGAPMw8
vncC5TOa9XRF+uyYty7lNeaEOia5ydbZ7lmeqLoHiWovjq3uN8fdZ1PD2XLorYy/
dW1QC3yw7ggRgI5afW4C0fxrUJhH+hr1GlilGxnZBFr9JdxCKTkduPSjB5mHtkA4
yhi/ZIOACFo8S/ihgWMmEhYPwTjDzKSuqaZxUr6XQ9JDSWF2pYBQMkYWztz5ALKK
HpqobmX6SItAbaBiBg33MTiHXJya/cw6zUHrrDLy4yIgXIZh+WVc0WBGJeufVxIT
flN05oSnM598Vx5XtODFEYj04n2hGIZcHB1A6CCcIKuKzKqcgRPRG22a+Upg+/a3
NL1AJpc1N0SnKM0cAChqV6qdNZx7VwYxf/rqAmH5SS2SV9wBDUmFUdIUzcGkAS+S
KYl6j06cMxyuxvqaE1wlNu6YPlh8vtgUBKes4P8uUTug8GI1E2cn57vco+aq/VEg
FSNk2I0zlZIuOOgEsDHM/ogS2P8GjSlaYepb1pmorYDF8XqbxaVOlxVPv80Dbi35
7R6cEg8x814+AsvaMRWknCJETp3TaVvrPsQ7fT9yA6zNuAehNY3+t5JcxXigH7b0
47Yc3DSDFu1Zh0RUvc/dGskkdh52nnuK0OehqQ63zw4efSdB5+2iixVOoHULOpbn
eyHJgPfIHB4Xj7ye6e/2yO3ZmMAJw4MalExm7qPkn9gj2AN3iZHjuK8D47YZjFKr
gY7Pa8nrBYpl3fi2o2r0w1I4zYEqfM2el1q2YGh+rZuXpiAJgCV/3Js3mzdrFPRf
4WqMIsg72w2B/LcX4fttcdWOcpAss+mFRJAx1GmrZlB1BEq2UzT1EvBKZGscByQO
dtBv5gf9buFHC4zpi5tLn051E2FF6sZdqHXHsYhLIFzlh2wdRnvBgSSqfTRaihuX
0Bj6FtRgorzWoi40IXaYtm2gGq/nQwkfGvDkA/Vj/9tle6LdCapFJ7KoASo8jebX
vCoUkip303Fq36ICNDuW+C8TdC9W74T6qErRRJJXEhprjJ63PTfimRk5xbnKwzsK
WJDWsCaDbeaPIa1Z3CpyAw3H8HlTGv34uFT0IJp6Ay6Sv0CIX5sA1p74uKcxwvGp
oeFrYwLPgEN+oyUs0b+KOUDtVgkM0mVQA+A3xPWMIs/x0lHAA1/DvvKy6EmXTksf
mbp5fSTK64h9Z4+Ek9aUT82lBfggpCw0mQoXoCaoJNJsGFvkmJ4GjdEMOrtVgpEq
ub2xL+uZxJr8jUULWMBURRjwshec2gaGsvVlghy1oCMGB17DY2qi0Wl7RvyOeL6i
duf7uYyS+k+mYZYKEya4XqzI6OVWW3Ux+3Skpu7ypNXPJEyLYVvfe9FDyZE1JMph
PJJY8M5ppGd6nrHaKyorOhCgny6+efAZClVzymn+PYwpBpD52Lifqk4ldNdTqXlk
t5fKfiejasVZFgt04VLnrpSgL+meT/roNhQlUcD9FwdZ8VNdoU47VYLCKfvBn7l3
uloBcx+1uNxeo/KVNgLP8tLlraSZ21mXyhTLp5kTC0rw9AKMoqcvSd/QK0qSjExs
+1QwBvKj/JehmOmpCGAx93mAQxE3BWGWTjmQYxs8aG8/iXzRHtf+xUcm3j8H0Ckm
ny4diYuB9SxkdJFqjz5r8Suaw7TZxV15KJCWsfwmEjYqJT/RqcVQWJsU8jh0HUqU
sCoa3j2bf77WBA+YNVopLFMWBAe5+q+z1ZT6aJdjuDNKPFTljtXQD4Kwy/AjjJc0
sJl9EZa/Udsr3iMsUvgr8wgdFOv04Rd7DamZnFWyPxzQPvZUgDwBrN/7IMXHVWry
1vEiZUo4Lg6taAhVEtOnKJxfMh6al8RCX7KykAna2v/I9KtKIW9yriVOO9wKlobM
gWNTYMoKHgRpOXaTfy4iHN4Iwg1mBsEmaHpfEwNAP7ZSMfDny0SPAZ6n2kmp3S+1
UuQ7fWM+KrmeD9JL312s6j+Urfpp0v0eMx5Bm1c+c8JiPEy8Qzf3p9cbqAGs7zk3
sohOUlUYlO9vVoHWae1N2xVNQj7v4CXrRcVYhd6EelwRpkKKsP59KppN72V8Mbxo
VxfNc5JsdeuDYB/xqZkkjAz9ZnVJo/LZAqf2+ZUunPQ7A5GjRPN7/0jMXY8EhCDo
v76i/UkypZLmHKEgqpecbAbOwn3vAgTydEzrmmcjcgMMO0meSF9aGz+0IqYcBAoA
r/zMBxlR6Ptk3EvnoT36pTJk3VV610LqUKNPs2/dOT9kYhHTaGK4MjSLx3YRgHDL
P2XdQUf/Ouo2Al4EfP+WXDVLV1JzgaRJ0mZx08O/o++KmWyh00OW6Y6lJqCUtswf
XOITQDuN4GDdJdHrkpe0t/+BlSrR6kitYRiILcJDCKXNVNN553fXQmNsqN52j4X6
1eU2kLtcJqDVPmKWwGroxoFpZrhqyEfqnBI2DqRRJOKdB14pi7HpDe/wbJTsQj7n
Qyeq4h4gAjHyUe2uu0e2xybjl2AmCQ50iZuHwbL9e/HI1zpjtREyO6kzQ7Vph6kg
EWSRzlfSUslFZSSU8/QzBHOZDHj6F/uCxbuAlJ57DvxTzsVfakC2O/sYemAgG+vi
JJxneek5dOP4go2FdeetvbPhpaRcTyutg15thN5TNTTlO0j56It6ml0DXDBzfj5T
G9i+O4OgEkH/dUGHh0OXP93ShB249xyZTcy0V0LZ042peAHS9I0cI8i33jvR4fZ4
U9sfPxj7AW7/MqfJMRoTN+he6+qEOIiEY0a1qCBV1PijeKA/FTcX8EkNPXxCg5yG
gS1Z7d+0z//024SeYgtZBjvffrAOnbsfzHygdZ0s/QFkg10ALXQX1CGpSSlnLxGG
Z8t//QoDVhVq2FSl7oFMWSxzpfnzCTUluf+5EO2FkYryTEE0ZxEumQ27VPloV+VG
YRu6POni12RmXh79SIu3mlPyfevgorZiKy0czMr4DhaXlc4UNkATIiPwsBx0rOxm
PB30BTsDk+0KQNQqyxRMJUN2HFesmziyrHt7ci08BG4HYxcx+Gvc0diCLoVsb/TB
Yw0hGV4xZBrUZfw16o4Ry9gn3RPm75Cv9c5SkpIEF3292Cm+Q87UPm5rP1azEYJc
JsIy7h3vmEUX6JPMAuFTPUuUnmOFStNzQxtjpknyMLRVRaO7tjKCwfRTAdDQBkLX
a4jKHJqK0pp3Gk/HVxHvxUZToso4MJBEweVVPdxQt6/UYN1DxL7DHrLgaNllb485
wOyWMT8WLPo7KNRBA1hZMFO6c1j1p00RYlWQQroofj/IqJtAO5q4G/qz2E+uhQji
o+lQZVxxS48RAcvt7r2ReV0OaDfu+yANDbd3iSTegp2OO+LhJkxu/WXTxQgJqtnv
D6N1hTDJECd0FsOXfWUPeCJVgj/+l1qn9vWA0BBRUGnGWbSYEu87shVFloXtttvq
ICj1NDVMaxqk1XLiVVjklEfUf1xlqIKIrG5Y97q17CJqS3bNXROHw7inVHc2f8bl
jw7j7U4illqMeQ1suSeRvtNZTnFVE6aP4xWLrC5QYc788BpOmJ5ptQfsw/KIHVan
ir8QJU9uHii70Rm4iX+4Fe7/TO2eefnrL7AXj/wQfI9/fVxJZr9xRg3TCSO+GJ+w
xtItBhPSl9X6EnSq6s60t9q+S7aGaY6e3hHsDaj5QMZdoNlhuVajbA6V/EOet151
DWpJCzejHfEaSdIus6EU2b6xJZZFnPYsuOer5G+v9oWNYnt2hvpskeEbjfevKITn
2m8evwWmuIQGpi7eA1rdPl5AyRhCwaDeTBe1T5MOa97ZrEgzXYfjOeIs2QNDdNRC
RPfBZr5z8IhwEE90cmBeNZj4viKlSPcc6o8kfCVdu+t3gXle6CSm7r0Jn0wbMiSE
3a8ut7kWajfRSJ4bZ8plfrvfJgCyLGh9K7Uo4UKLFD2e7ZcUgpB8NzhrhBhI7EAc
xLi3SZnForjLOv0aYI92UkXKmpxp+ivtlIDX7/qijsIJKUrj92GtGdAIHa/hX3dW
HpbqQ0q97eoGj/F4nxLY1eiLlXPdNT+0W9NasPhq4btUQWw6LVZKMSBhGY04MBdS
P7go9U6+UX6Op9NS6rhYx/Z98wGK/gmv6+CvzaU3jPIxWpOfMjNZIAYPrs0ibLLW
/a3WElLsPca02l6hqqCeXMTadWGWVRM+sWn4csXCv3bRIJ3T0INMZ4nJ2uHFLF3p
wpqCtjpY9TePvSQahTVUYuzTbOgMLvZTb4u6ApLnHO4HsRuHhWGXF+rb6p/LKNAU
SuVl9P5KU06plSOsQQiKBQs9hFkkgmYSL9ZUNN85xeZhy0b3xq6wWoJiPWjXkWzM
WtqGeaCCj4LbdoLxtKhjTN/AJfuYMTzixrNRISddmeT5Kb0/VIgqUNg2FcWvf4ZJ
q+Xb28bFLfGeMv0GDdK6MFnGc6rYvCZaH3W4GC9j2IjYT1CKgDshGvtEZTd/7boX
63HaUS6zjMtLhaZ02TpDodjkM11jQecTkB6Rq4yvrGscrqi/kvHwgrggnaThhAvW
IfRfYCKcdKXB+//fguYa1rpiwhCxbj0vQlRY6Zb5LCXPEdn8MYa3jyL0FL9l/Jca
nvLq+yd7W/d+CR51XG3ETg4zI34VIJYl5r/pXiWrdxu85OwvS7pgIeJ27KobO6OX
ECps/qAw9bp1J1jCZar4p2956I0okvJsdOZH1RfXOGd5vI8HyGlj+4m8ki/sMuyM
3SofzkgkL/KthGq33g5e+3c81xcivES/v5gCgN83YVHUKOCZciK75yaYO25EC4ip
KWIz/aLQnJccfvb4EAb05Z7RBOKJrQhAs1fb+DwY4lIdctf8gygT7fnaUWYRTJFe
O6Hq1+J8qsqbRFHwnIp3RJlrJFuz9JDnWLzv2wMQ7ZLAKp7FeBYkgvGhMs7Fs7ff
sta1Btc5LOPatA9/OoKObBd9PPrf4O/2pOCa5clye0zIhS+eCzuzovrrcYe02LIe
Zn1xwCvqOzRcIGGBR5eJnWTj5K+7HK3+7ULctbVIauXFVufpdUOIxXF+z67Agqq/
Z+kGoUzZNMBvMAq+v8Vx46uXf0i9WMwVV9AhRkzFDkD1+jlU0kuK4k40V87VuGGT
gsln5vWhzK7tiP291Pmac1PLbW8G4Um/kIREJfG9tgmI3/5wY81+E/vxkn0B8w5A
2Lh1SBO9xSg5AQuCo6B0GfIjwtbWaBSz02j4bqt9+IkcRhO0FOj2b5HHYL3/7cOq
XjnrKkiR8REjwAJBA2XJqJKHLlLBYd6I0xIJZeNfnsraXqyyTa/NZBkWkiN27zbT
RwTkSkKp3O+zcXrtqClDYqSERIlPfi58OwoJS7ezyoDn+DkWbNIBQy1Opx8ORzvE
ivO/OIEajPjD2eYsAyoCOMgJH+rf3y6JY/6kl3ukZiTN1KvdtWvoa30zThP5H9r4
ZtF847gXv3BdKVsgYNGZmkPbc7f0jqBUmxVcU75om/AePlDnMfvYv1nz6JbHlX8X
e4w2rmB/2SAEKtDgDWsNM/4hucSdquM08F71/UHNmNWEXBIMibXZ9LnoPD1aPkZr
FGxbIH70WgBbs0sOyVIemO9GVBuV7FZUSJjemGVYE7fNxwuxec7MvkE8e5qP6b+b
s7dtoFIGurESRAB5tfehDY8Gv+hyc/CN1dyt10ymm5IPYwF+c+PYWaS7pHuVYTOy
SG76KK7rAIFihrqYRNiNJlqG91xLwwMqW1OAtYjMOPeRvKvkLvfQTXfqAtQYcUwO
undigl9DsIbfw2CgkSA3CuUMqgCRPOXEQlP5e49O+I3FLeZkrxqQ4BhVd9J+eOk/
P/iSekhLMlRK3RTfLbadaLXhWCFtzee+hdsbBEekL9qbEIT3J/z0kAp9yeW8lhBd
3V4J+soR4jQKEeoriINXLce5nWKIx1rOpHaB2icc9b7hKxycdtSf684BVuO2PMaa
t3Hi6w2c5AQvrBw+k6roBwnkYDUcSHKvT+EuAOOCUsu0ILuZahtLFeFPqwjSwyEH
TKz8mWjyJa+AkBiTocV5Y83D6P7cXKgmjlrxqcERHkMYzRFto64orbq8DWVUjsyR
/XWrJyuuqhCTshykGnhboO/Hf43R1axpz7Dw3mWOeHUCBn2eqRULeNfG9i74plqM
5hxg4AQZ1IammsoWOaLAwk/wEmh1+DMDW9cC70OhUTey4UuAkAxSAA4ifpANOZPE
rrBXbCtz01X169znb7IMbkdzLoXTE1t8cz34MMmz4aJurC4HKcL2i9QHrwL4BstE
Fn3c165LAIHYaMmfWRKuhKSgyFR6Sp6YdEoSXTNm84+Y+myY98ZZLmHHMyJ4tHRf
GQW7nmalFgPF9viGg4zPIIWe0nkFGQOSMghrvfOstVP9B/CRZrXJ0qar8HySkk08
Ja8bls3m46yIRmuhn8WE560zLhHHh5fBQVLnCR3JCkn0ohpxRA9TcgnH0nlyXv5r
1gIln4L9XUqYlUI7n8gyhrA3hqDQMlMJofqJdT7jLUD6PvgQ+fXpWVA4/1YtJnNk
ulTfY/PUgW2GTybVPNBodFkU7ovkBFyCBKVl2eJrM+SVWzlhPdA+yJllTfVQV1b0
871lQBPpiVNwUdOEBj1L9I/4iaBEOThKgc8dwhW2NozSRbXszh3GDjGnU6eXta8Y
igHSPgNjBBVv8hvoCsBH1nXIJ+enCJvF+6XnMkEUONjNVJsKxZzy0B+ULuAw3+l+
S7XIJkrXR97/ptCedHQLwBbFJiHmZ1tf7a6Yx3Cj7SrmcuvWmzJWUiJxQ1rJFxum
rPBHmm8K0l3M8qqukDw9ffdO0tsFxgUVrGZjnE+RarBecQ11snZ0D7tojI3m8yp0
kN7+zlWiEUsaYNpTV7YRvY65y6eYHbM3zwoIfWFp52x9dOEGdqKg6Gqt+BjluGpJ
Nj6R/bXqbpBPQwBN+/h8gmKZI3kGlUd4spvmWS9+SChwa/SGrR6Dx3eb2Y1TWRYW
UoyyZG1av/+xO2mYeK3I53PdI/2x2VM3yDvfC6jWGimxZ0oXmHUNo3DkJS0qBZtP
FPwYx3wRvU+DlXUVPoAqiKRghatGsJLT0z3u39GR8pgrnF0HqVqyKfKvyJn77B24
UlHGZz2cGFhaVOyETWtbfw1KCUHNQr1TOg4/CSYkmnxjJBmogF5smaRB9iS8OwBE
MwOHBNbYgCAHsmxKboXM3tFPtdSPkHWqNq3J3XEKuFxwjr14OPG326tY1eZjlj1X
UyRvLlCt56FdJKNnjN62HqGQ91afXOooSIP43u4HkG+sgu71f98vFpODnIFcJLZ+
EjfAgoe42QHf5LLxmhpp9P9h5etVQ9qQAr2ymZP5sFf2La/JttgdZm4R8I1/1vPf
K3Zw5VIQJqsXyX41dBg5WWKZYxQ7pizRAKPJ7kaE8QNGMVPHSHrntUjBWsYSGR7l
69AnVem5lqAqgzVKsarMFUuIp6UUkOwzxUWWEHjUWVS+TxNuONO9RQWaIqCG8WxI
225pympDrY19vs0AL5a6/3tirxGrywnbuOaQ6buxi0GqATZoCv9f38hEB1GYUy1u
pdhD0w9dNKFZn6Hr47H2gU07Po7brIHf2URpuIRpV09IZPpGsLE4OKSNfPiWIvFx
WRhQfL1jWviobGbI6lhFFFwrllHsvwa7Xv6nkKYjfB+yu8E2yvdDseTayKMU31UO
VwfAcEokrZEmmnyzmomB0VO34yfjTZGTfnxX2rhLBrsh1akaj7A8RnQRHnvdXsXe
+Nd01eW+9igq4W0sw4qAIrmpq/s7hYiyNZHzw0HonBClmSARCHJM9/SsYSMkWE8g
6TI2FW4uI8a44b3LFQakTBwAphsNms3vy+6Nm+/1XgH+jBHYDz/cOKSzt03yjw6e
7utQVSRM9SAmTBfkBFaGi5ovIzfBT50D1+iRiU6iMyS8vnx405x1mbH8zmDUXKVI
FSKeUpl1q7OPPyNMO5aERF5fZIHTLfZwH0t8yHFE3EZvRxAHf9p9e7sUFMEorJO6
PrA6U741hRQNp50u0RTK/h3KECTDfR60ZDtorscL3AyZ6+okYBVrGNvRw9dAJ267
R9XaQWRqw8r1A+zmuEBQc7Ja/Y80DYPMRo/s+kc23tf5kePjdSIwmQ/fBPuf5rEK
NiHcmso8aHfWxLX4Nikl+mrD3jKQtl1KSR6Iik3zKrht5lht6jWr4Em22yfuoHVg
c7tVBPQbuPG/grgxzqpc4RvZQK1gkg1mMM3vKrWcc7REJv5y6Kmr3rSKSEMISN1L
6zrNGftlfcs5QO95m7TpZNjLFhiq3EH18Dc4W4iYPZ7ZDj4tO00McthJ/CiGPs5I
thsM09OmLIpfaiVhVDOebtbull/mXJHxXXTXmkFkOO9XkztLluAv33i9rPWq51OX
ZNqORNOALgxpghtogyJv7C68FwceITcI7fG3FlK8i3jaCDTSOEvoPTw+oTX5m38/
y/5a9e8KaSje0FpDgVqwoDBPfoKTznNkhxnPY+iJ6L08fIdkSiLPrPj16cRULp2n
ZgFtrvPKI/lpzJLGFBC/iBHvpkA+calqYil6TmCgp0dwAmpzZ6eYlLfjkfGC9VJy
W7z1pidACNHEgsoga8Zv56o9+TcnV2FBOCvu4ikq3gYsLXrN+8P2y+AuqVtxmSL5
Cxu388ykel7NeD/Etfu7xlbyIOFif7w3pOrQtGIbMWLZlvKMgtZzF1pkGvQduSgZ
D0tqaZQHzExaIdDrHCtKJWYHCyHuMMoc+NfdwXUveuyZ7ud5VqfpIOUBG2x0+w8G
+H1Y7TzFOyyNnr63wJzbOWf2e3HlhoI5p5lPKMItTrCFTI796cYSDIB+LSmUprco
5iYILm4/eMGa3pl28SjY6vNBiGy1oGmTjGPlBt16UNJ+hVRtOlRomATatN6Ul1yS
dREWU9WlzqtzX07fyPZ9rgzasi9BYwerMF08HMrVBJ1+IGuBuHD/irLTbPfCBYlZ
A2IwZQWmPFEy08VuGfVSpCdUPmto080if9RhRCLq/csmdgqMi41IJdr9AsnXkv4z
ClchCSK1c6tKx7JhVin4O1xDxnbAsn7q+ZiqumdxOWlNzI7FZDXmwVfCyB9hqlLw
R+YjU3h0cia1k/FPCH/rb4mGdk3GizK7r7fEO+0uuem5oR5J++/BO+gh7aXWX/ne
30Rphp05PyV/HR0H4djB8p1zcyOr20MGrGvuxWRXxThZg+i+qn+mKgYSZygue9qF
OcxuIaIBUw8LqySnP71Ss5Zs4sedvuA87vxgSQdQhquJorLdU0Du/z9d3IelLxnC
TZ8Ew4NbEvsOEjfLEWCBOzH42E/W91dWZQstn0AylfhHtlBoaJJfjLla7+osPzB6
IWMIeCV+y5dp2stYosu3QCPRO5OldRUjeUDuCT1qp9Ko3tRVRObksng2j2MMW29v
rFMHHhFc89IKgE7UhjxU+vkiscU2xQBTPyP8r9jf1LE2+nrGbJ3i5E8QEpawqPZ7
Pn5LtyC1W2fJq4Sm9cjF4UlEHZoG7utTQecdD4WHnhGaP+YNyWFhBy+1zV8FaLUL
EHug3Bxed9EdfcZe7+HJN2SgY+CDOdK65b6eV685XhB/hEEhxtkxcnTw87TZVb4L
9d0cWm7LTB4gHVukhHY+4iy845ibrv53YVpicebihGFKvx41qu9ddXa89MC73uNS
fpn2nGgCR40xRqc1q5N1o+5dv0ijATmX25Omf+INraij4dKy0S9AsQOuGSlcmwzG
YuY+h7ze8vBAqK2/xeyRxodN9WAS3eyZQO1itNoBJeUsrp5zSHxiK2Ox2nfVN0LH
h+K7Rim+zHVJ7LJNhygwMttvN28Jj9fWZe9nOoKR1c2u89iJWY9XjkLKLnVvL4xz
aGXwrA3veL6ZrdYzEeJucpLDOtAJ+S4/wHe3IuVtuACsKnG427nWNSQX/SG3KeOC
3msuWHpetYs9xNJgDk27Z+E4eczs3FEUKkarCJVhOmtfnt3SYVGhXhtcdddmaw9J
flOhzGdOfm06/cB/AWywhMit8Ek/jfaxXCqnDuzyfwtuoUSO1m6hePMNGB0pwEAV
qbNi25GFNhjCdrvIO4nlYgegd4bpGwaxlgGUhcGecOSPCcFKBObH4Kisdk9Ilq+9
2UwDX+jtuNuIcfrXz0825a/jAweof0otVbuiQgEfMSdt30P8KhL5uWm72Md9supx
5ltIfIBKAFrd8qOYsjZAWSsG49CkVuIdNPb+vU9U2FwS6m01cJHw4trz3gYKoujt
Q94Ecx+9rHh5wdgC30zqXsVN05gDWFkkS2OZh0KHF9mO3gACnq3GjPst1CPPZ2PS
8uZcckC2mY/VqOiem2tnC2rE7L/junSi2eUMyikoBMrnmoGemQKU/Oi5j+YzIkOF
OjTF2bAVFJUyPuGoVCC/7+yQU6pcgvjgpvRH7p7ZQ27y+jHMaNNflpc5zvR8PSuZ
S830tp9hI2Jli3c+d8Db8eomozZ99kDnIKe4I1L1llL/ri3i0lIwj+sMe+PfRWnA
6jNvQrtVq/Z/Ch8LGueve4BorsE3/oCqb4Xj/hhpHP2qAMcKfZM0OUq8ZvkrlFNY
1QwOP75q8VMfI92MayYnjwBexhIoXWxMpBbXTtL751E+55qiM5HRoHBpnP80buPp
mdW/SjvGaOtRx05ykqhXZ+QRrr4JuLVvJlEi07iBu0GIiPbe+ccgJp2KwAprG9Hh
Ax3+4qLcCgDjDVvYM7W0YIAbS5nqRPcXRjcHavh/7Ao2JBgzpnAvZ+D2Jw3NKB0h
jIeNXdCkAJqmnkCMjC3VHMtiqgVNSO8w2oDuQ6MyOZno9bOEV7tHx+tu8KVPNQZs
yDdURxR0rTeSJV+x+XoddjVPuGo9id/s489aFoTABw2Xv2fgHcAFbgqGZypgu4JC
HjKox904Gd0HFCVJWuORK5C7sL+IvA5BKqgaNXgeyOE/kO1O1WbXi8HGiNCEkKA0
PMWAtWydQRSDZlUEiww6EpMiJxbkNNyyZGPkhW/KeWIXmbp9KJ72lDkbE9r8Ix2k
IHamlO0xnSYaB2Z8Lw/FBDJmjudEq/tBzSPm82BV58WaYftddvs+7a0HScwo3n31
rdc7PHpRWn5Pk6mRx/fXNTsS/I/0pfpuRTte5jyeVGz2iVCWNRjbX1GCDSJzR6bF
m1QNEL8TWJRdl5TFnXtgXZsG2rgxCflbYAG8Q3i5P0tMhw+Mgj3N7Prrc+ypKt5n
uHTkVn5g2a8A5gOYN8wi/9Zw38lrHv8Tnn8Zz9b11/thRyPtRLAgI20dI+r3W0ps
oRFuKVlYdqmWrfau81N3ZDJxpFOP2qdYCUm86G91MxE8BRVuVvL+DgUZOmDwYsid
iKQAPzz1OWcmEDzVCbUnHxMBPEMNIbkz/yrR6MTVfIkYuL7jkz3nAGsOWc7oROLd
FPIrSzQGKGqDajyoYtDfNZEHuqmDdJgQtMdl8kAexBHwTUjWs/UwEFKmm8Ayd0jy
iBfnGlvy6DwBHuigJDW8EvfKPNJIgEF8pGT2IidPLUntRym+f4nC9SBsn0xad2kd
oXdGG+zOnA5ZlLk/vYS/bNs78TXPSgvLA+qflr8pnlEzSlU+xt9iOu3hHpHBw9Gy
pZz6HnfmiKNT4efHeJpkEMSP43qT3BxGtLiQeEV1Znx3OBoiC3KiqGNvx1+3lJur
ZkTuFlmvSh3ea0rjqLHB/6N3JUYDOTXJKsziEgzDrYPazw4qHDXtPj+AjBBZkTBi
24d/vFhgyWZP6aLG4krkS41Ex1dp/dr4iEn8OW72ZwKHJwH2cKWMn+YWLiWQdEM+
c8Mru8ZblgJqvhT2xjWHRoRILxOWZ9VdXXyX2ZwDhau+h53snPm3a9//NFsupig/
E+18xb4CL2tpcVAZmqx0s5E46sBvzwPAcKzCcolrfvxErQTqyy4c3g+w6HGLFYWx
iXt54cKC1BUMrHntLmPSFkDdnsxPkOagI+FL9CVaogtjOi+mCaUxnCTWsK8V+SHq
35DZIv7WJpzta/2QiJqi6PzxLGgijHMFN1jBRARBiR9X4qjoDLtACD4km9aV+uTa
J9xF495cG1tlqUrPXih1rgR9zCzdoxfbv7wVBBrA8SYOzum0j46Z6eP2M/lGgxBl
geXVSe5e6v/0y9j8taJWRu1Nu/Pc26yNRws9Ys0XFXDmpMbBSpr0Rkw5l8hT7WEA
+c32zHxCDctqy1optVPd1EqViqGcYFOe5WJ0Q5AxETN+YfdsQ6wFrghu3l1YLptM
Ew4Zif1ZZPqrNSZ1RIc+/9DGevEzrJyYL240LVX+BL220IRw0xCORN+35r6rwWRU
+cg+bxdgFnkty8lRwE693AAK5OS51FQaytXUtp/dmDibTmxnqjq6OicXRuGT/OdI
ON7fNS/pz2tTWKyIgjD4Cpv11T8aoTFrSIExB9zciRs6ceTyQ1+iybIER7u0CWLw
T7KMOogoFT4SClSVABF/b8cdIcprIR1dYAtVTCSfWpNE72Zine5LWWw8xiUM2meH
JuetJwnIiolwf1bYhtgsulwqA7ZzYpEPbzNZJ9uv6uAZOZT9czmKhoaUPXa1CZtT
+6HDEoQEjBmCzF7pK70M1GJyV5b9cz/scm4PfAh5nUEjb3xnpS+odxa65ixZnddj
rh7Ehtg+LIpyAOgLe2LdNm3rBGTju9MuZIc49FR0jE4lSyUuy3YBDM3QvvCbhXYl
TNdqKuN+Ub8x6DVjyZQP5dXWOt1DUXVb1XegWF6fvGAGUcN/tckTBRnNr14Cjlg2
zTvcVTHAH8cMV7z1ff3Sj8GC4uCmHNbOJbO9yIQT2mTTC38B+kVNmfk2vxgMMboC
HCHGDe1PF6ydyGJnioveEc99dgZ72cb3HZSi1S78dioZuds8jSf3MafX4uLjOObx
Maxn5JJPikyHeWDtUyqMI7b6rUL3QdNp4PGivLzcGX+VRpb/kYl6RwcECb8DrLd/
MKTOjyDwPE6DzK25jWBeljG6ZIkY5xEWhCp1qyir3B3bVXdFKYM1IJH/lKEtlB+P
ApHnru+F71YwdSJiRVnU3QnbAIOEeLGdgq3cXtnH3FHu/e0ixDbtetBqIolI2dnd
rh6fhUvFmxBVWosKi1zxWUqgcJqVTsooha80WVlxCcX43XZRXrXPmH/C8qz+oH/R
YeJYfneDEMBNXM9uwFsZG0ww+ZCp/NO8mZJqDStYT9yi653Toz8oa93pwx4m8fPG
1sfqmPySxZ76QsgLMU/h/zwiZGzEyay7vXs6epZOFHQUI/bwlywzdKgJTxro+TAe
Ufd0TewduZ+oItQTentCam5RjC0odZOVzDKbpWR4vhEFf7HPIdzdIuP7ccfzvu79
UefY83wabmSPGe2rrBfSWE/KYqbF30qoPjsnCiT+13Qc9+eVEOeRQ2mf/GeLDzxp
cjv68lm9osPxpP6jCe5TLvrFpzWsGd+1Dnbvpj0apEkchXR/8f+Q3ID36GFCOIrR
cCTaSuw5OWCfldEK4+zzAu9gQIX750RGb93snDumv4XUYM39zidx/TBtRYYBuRnZ
5CI8sdcalAiAMonkx7BZNNmDYi2hGIAY/J9b33DvEJZFRtB3jxNr1SGH6qSTWWnC
B5a7HhYtEIM/6iJF6AcoxLOUHP+Ni6vn+WVeDg5xm2lnIXaEbivWz/12YD77Gp/+
WDF9pD6tkP5rdTrh2QEj8cXniSlx8UE4xD5Z14fn9bsbY599pZ5Es32Vc+mSILaR
kRWe1F5YMz/l+SGOenbMwjsHTbchzfDp1fNa6HR5iFAlTcGCTVjhL8e7lX6UcK+M
/3g9S1V7S5Gy2A/snEtgsRmhdBSC3bh1V0H4KoEyalFBfcmyCxHxWyW27DFLdRcd
Ve/Who4R+sj335MKpB//1sru4LOvryUVOUM5jCUrRdBN/00M+mMhUfhvsCQBogfK
Bc49Q3L5cq8n0ArH6id9SGVU0iE/cPlOB80CGujL/wkPxzhEo3xj8jS25bY7Bvrm
CLuudoaf5FWe6khTm6lDwtISRI2QbRhdIxtVNfChWosW0OQKKH4KGKK6QNUbRORv
5X4tX02SO+wtgKj2qAn2bD6WO8WZsOqamz8JKIEw46tzRvzO/8ays90Isa4faZY8
EUl/eN2KSlAgW4wLyOyfaVOhPEGjqnwiLQD82iqUGgmsMHmUmGWjWTCFw2qylCML
HkmvJbngGlcZ/AaggFdMvxGq0QmQRUR1gag64yqD3ScwRBgUe1hvRQBE3hWeWXDz
gss1ryb58UkrOOiB2GREz8/pfw1apkFbhaC7eaFTex6nGGCI8+sl256X1S+mPjC5
ietR1s7RKssC4N2QknrrjnEDr3bBASAV3A1SR+ge236wlkWSZjq2ujiTByZy8fGf
YMemD9tEVZ5ND0LIKwQ/dxE2jSwOsRoTHcWHFImhqtlNu8ONkGOiQfrbKbZbKuqO
tI+8spInVqFAdwKNOWeiSt5KaVmSZ4vxVRa0t9JG1dv9wJnIGmawmqNPo2sTy0JB
vTVhyyLudg6Fut4ngIIKbbmYlm2lwM5iZrXSVNYs+ji7aGrkMdFnrY3AyTFA+Dzs
dx6bYVd0sqM+RVTcg9C1e17cBPrpss4rnyaCBzElvECHSS06KZEJGHfQZcqoHMaa
e9AQVJ98+YZLR/7TfZ3WOr9kfERPWph0kPfK7DGyuSC6N0TGgrbAHgpsaTYkryzf
C8iFWdAUaxBBg5A+DzqLEPjrt5qUOBkE3WVFGan+1NXQZywdPlHxkgWpFFixrSoe
rEKEucHhWc83arlB5Koj0EQKVMw5fRW49TQ1pTOHB4wB3jag0D9QYsIYOCBGu5aG
uxdEcgBaJGyvZgsEzCyUk0n8sdLecO3QlNnsyNHiWgIlS0oIbO2eNAAs5Md+7iv9
hr1f7Wif5579bFmC3w/sidYza/kCrOVpEsWggpo/0E72Cc90CN3YfI1WA5JAphAo
wUwozSrUJJNCfoT7mcpdGjnfJ2HrAzaBf0eFLenYnlA5LKlWKn1PoiJLmJVOLEC2
wg3Ngru/XItu4lPuu6ctKS0e6dkPdkkArG6+9dngIP2JDC4O5ki4lbkdXDbi9BGs
Y+DjzwYUAvT9ojLQ32tyoVpIUqPJqPiO2tS9jhdU47lfbAKOeYlS2rhhEdA9azfP
5GhR5E6DE7cQAZfjoeiz8/NXO5qVmpst0KFO7kuEoxWGyOtH2frkptKI2B1hSip7
sCaB6QEAxgyh62TIN4m0IuD1mAU9EcB1Lv1RpizvvoibewviCr9hvkzEEDw+6bNT
dqFJ2tlcCn8FvCiAunL1h14g03rARAKn4NYrxZguDCsIZL7adzKox61G5MGPGrIl
+cWpxgh+R4Gp/wyxPGwzlIGD7G/SH25NdR0adeFneVhXylEz2PWsmkyImcvyFmFE
6JX1bvbZ+VmfjNRhde2N3JLJ+po/kT0F69RZhxwRW9ttwwE+hC0iLGM84205uL/U
BoVoOPrc98kBtopKcBcqkz1oxJPgbsPlUb7vUzZSgKqLcUPcPApbcOHxzo8bx+Pj
IxjyDhNG4xJHohu5oN8LZBeira2y0ypubDrBs81fS8lc+QNFLcxU0X/PGkxryfRf
bXllp+asFf4y6TxpUEMzNKoBLz0Fz+3aTB5UG+zcawzvA8owSBZc8mapPwMTdkBC
jFpMvfe0W973KwVgBy9qZspFvuivfreVOmmeVjNCiru3RjNgOdGseGe85htCtd3v
ijstXwTPjQ0Vk9t1kKBo1iHAvZFTVnvq6sDqSVxhzNmp3TWIxjA8BKOCB9qB+Vro
nqY/V+75UABuz+94rNVz41xEMwLN/Yd0M0oDhuzT1auL3pYHksafJdQKpL6csKrY
CN/D0sH7D4lvxciDzWD9jTEN0ZhEOaSvStCOYFQ1ItKqKg1lqnoEdBygkcNz5+WR
fEY1D+hlZyc5h4UBqSkUQeCP4jdv0KqolTBwOem/FiyMIiDlQWtMyun7yA5Y9jS8
Sq2hcAWrQadSJ/HRfmVVZVXTn5IyaI7q5cVos3/y1VCaYPUg1Y99sUuJiWhdeV9k
+bbchsnR5EtShF7PpIBHrzfGpgzQZhXIZOKfX7Ibko14MYbHEbc6zi1taQtGw2Gn
RoobKGOL/N90mKNGr28et15BtRyaIHdh54oCialNWcB8cNVaZaEpeqSxHS4HE5Yi
PFFlGJvI83hXoQfEVrDG0/rQzIQt5EoE67U0qr1vppXseLLQik2smsisRZSgIYbz
f6KpF9WXBZhuoP/INcIdf1eteMSWc5xRnAfNpCFWNjhUmG8AqE3QKj8/sS283nWg
hltl07KsYl4dSORhvU5pOd0LXYgvTgNbtrk6eScl6ww4VnFyrcSZ4e3NRjfDuET3
Y/QEX7xhCpC2cmCtvPjOK0TRyX0R9881cwvqrG84Hp3Fzqa1kJDdzQkdP/eM2onk
LdMVzDZETqHGu3XHKO9LSDwBc8L0NnE/Xt5pwIWQF1Z2NOsHkcYksVGf6cRQcu4D
wJcpdJykQwMLUbwecNTt/9plV2N7X6Y5fIWZ+FNBrhTLsoki8xvMh9eO+OA0hfQU
2/h+6B1T7I9WpLzhhLKlcMM4TtBYximuVgxwgB51q95nTgFGGUbXQ44E/Ppb8Mn8
+TRX/WU0NpQV+7K/kZYk05lt93DX141oL1A0bYFyLS2B07gre06CZBy26mJaqjqt
BF1pViQUg3ht8spv3xmszO9Fjm+F8KlVdHAufgo0rTUSuU26gAdKZPfpWwVAm3Je
27sNlx16Eg2qEddqGX8I0sghuUSm5XPTJCm+7e6OAk8KX5r/r/Ts6fW8/3UXj74F
+OTe8V26Xirz8ELvCPyRfVKEVYCEmCIsn1i4OJlxdPlTsDy9/ExCkMBdkscNLT2y
qlCJgL2qouBL5vGAxrsZeJKu7iQJOWVOESy0jGbVDf+HzVti4NEftlcipg52auXq
sVqjmJkUcyigZgNp1pAxsSKxk9kyEytLdELaMEfQS3jR9eMk8WBQetdNwl9w61kV
niwInc+Uh+lXAzqGGEuZxyZlQcc9GO9dm+IodY0cUqubbFCVgo/jgvzfHaRN9Ay/
n+wevpIVtHjNKI0Lx9tB7a4L5LzHnTN/ec1StaweRKjK5wvW4E+u6BHwDetVp5LM
qzK4o8nzK7msSOLKt37yYcshG034yRWAposI+04gbsjpnZAe7OcuR217SPwLHgNd
LAtbOBE2JpCZfllaw39DBe5nvMKABLLatjPSOI4ejky4irYs1/UFk6nxGSdVvDe7
clx8vyeSjDttME7fAB+KVcfr19zdbsUqS2fW5b5G+Xgagu5evkjU2Sg8Zj71IAfS
6dl59OAFYWYDcaey4ua6D1YfpFfWBNz5Jk7HdAlSIjpX6PywMiqnoTp5o48XvWqF
Ek0u2Qwa3vrTmbjEaTiKz+T54w1zle55j3B0rq8iE9eQlwtAWCzV3LZLRAY13eL2
cxgj3meBAwc+Dy9Yj5XAfNoJE5ZvNDYGIIth4ghEdLYSxSKtQOdld3dJHwcYxxFC
fFEsGFG2KfjPIjJUOCq5vMJxwsPhMG1XzWxHZat9O7yeJwF+tuNHXU5PgenaIcwS
5V7QYQkckTEvDDwNgxAKPiBIJQljvYC9GMIlaDgrwDUzO6FEJIWfj9iPWX5Vq5ye
gZ2yIiiLie2iR0Zz4duABtp8k3sz/sIJ0gczyp+KFifTc+8aayUUYoVedvVkQxug
v4VTGpje8/WytTjZ49uNfvln3jNI91SPCxRPijvWcOA1cpEKxz+RWissL2Tro3Ei
9EWXDsC7c9vx+L9eSpzbrzn90uDhgh9g/NVrH0f8P/THdq1kCcSlWYuQ9JhsaZdd
Ajn/1YQCAf3nWzy50ghf+bs51UuEcX0NLhbI5qzoM5/642eTbtpTArfQUAwBXf4G
izQM4XqQsv48QMnK0AxJr0y2tz1rAP5M3moNhdd1gMqDUuap+hsikCdnFpOwcut1
MbM5L0zD2zHa9B1AiNei5n3loEjVNrE3zU/FhUp1sAV2B+7LextR8+wcCayplbUl
VG9K/+2Dz6gXkvKF7b/7RDgwnHIhAz3jbO8SBcwHNV/CeMV9p2l9K7HvJAFbI1T7
NySTuSAbM52jywVEIasVeQwsVMaPshaH8K2MnYuJdGmNVaKzsWR8zShfdv0xvEtV
E30rBdNI+v7ugnPiWONIKVs710WWZ2rpb7q4NwURJFqRqa8KXmnPpRX/58tVVBMe
RUvSwAxWGVtL7rvXM/sE2uNYeVWBS5wmpOKWxVb4jdXVLuLoq1pegbyo66J0qTdi
QbYLYR/Q2U3cjjYtQaSCPYVhk9AXXqYnMY1cKyoXjG8Q7wOVoVjKg1qkKPBasHRF
vbJ8Wq5tm6aXcaq9GYWp1bn4UF6cqWP9Ky+4eizylfXqd3LgOqub+4PzzAMOIsMR
w+yJBGP+iX3XuJoWia+s8p+DRbFXZZSjG+FUOgR1l4lS4qrsl+tK+4AiImz/gN0p
67YbClSTuAVAPWWw7wzbzBMFB6644u7/2mVdr0UE/v0ALKjP3CYbE+myz9wVLO3o
/jecnmU9148l0T2ZIqsqalws5TiDJ5qcg02LN93yahU/vHYoPUl2DrAp50GbWnuH
seahzrLhFOVDlrZMCZf4LAe6f0v7+48NP9Zp5ZnGe1RpwvcMxTH834DmlgH42SpF
t1VFVBH19FTNMvZWaeqU11Sq1nZVy6DHMi8bpDI7KQeW/noOfVsXvkjR9uizghEK
+E/XounVz5igtUbrvWRV1XNcNQlZi214QxNHplw9Bw1vDi1VWWUgWEPZ9GPZ1Few
fn+tQlU4oGdUsmeno5e+cpfnAdpcPvNUTa1Dbg15JM9TioteSFXWG3Hfkrz19C1k
mwBwQf25bzyD5brZI3AVk8AHCQOGvLiec2GcL1ivR9Wu5cZbAyacWGJc+w14UKXs
+g6GURRbmC1uZCOX5V1eVy1ZKZxQ1/ywK5sbfXoAfuVLU/ZDoLcT1ZfwrY7i0nzV
cFC0zb0HwW3lQjqWPiBNq26kcWJ3pNfuX/geapYkGS3mk/tIpLm683bZMlfEcODD
NK6RZPgWftjc8WYkU2CfXjaVetHP856XmxxiU+yUFwiIlTuHFYETHv8m9/pu2sZ/
xJ4Nhlg3av6yU80lKgMnjzfkTQClU7NK0D1Gh2mdj0HruzPxHPrw7YpAmyOqddfo
y14qxTTPPyumyffgel3jODCj8ouZSnpI36c8xVlYGiQUUt9Gah3GyieUlVcsj+b6
IKFbbFYIJ9egZlCYhdMdUtK+gRBmgEej3xx/4AyHnr7eCEK+7XEcs9NyV2fKELh9
5oU9Aw4qbUwnVQ57Ads0G2rlgdS0BYgM2QVA5xfhcGpqHwd7tE+c1BV6VX63eR/2
xcWle/f0SvLxsVYkT9zmMLN97hVQ2qA6bFFqzOb6T+qi26nTMd4bl3x/dypBbbY0
sDVE/hZCuCvUXEKuEX2U0PiGdbdKx9QhfasJpneKQP9ZxmzjeQEz6UbpQs4IFa/7
B6pj8FJ9d2M8UBuWN3KHbfa1+EMqq4Lu0/7fOeP/3SiuMpaWEC74f6Z75mp7Azpy
vyHXXxWot3FDYm6vXlw0hav0bwonw/gltmm3GhkPVOukEJ8YrwOwcS88HOr/cM2u
Rn2IAf3Py/ga0Gve6QdAjvK9cnlOsUwwq0QSUe/PS6mbxPM8/9Sh/1NGGWihvFAM
0IW6/AphmPBmTGp/SOn7wnxCGth7hBYveqwdZicvs178NNJz/9aWnQNNcn16kOs4
9l4OjlFL9qlSbx+cGzpZP+JRtU1fO/R+/9aT7CJFETPcZ+79a3NsJBVdAgurK+RI
0oihuzUUw5OklpmqsLL3aTtpMWYyz6E+QCYIXGFImJesVTb6BF+X2vQ+8pgp88sm
5p/81EEEQB4iM76S6t4BbLpPmhGpyA6LmDW9aZZAbGZ3nL/ID8P6ppCJXgTpPcfr
EsQMubtPlJgE83GFtt6DO2G/eL56IYRrH8uWbfMymzM4C/9Drhqh8A1RZdXnMkg4
75iSCoQwRP78gcFVTWMqkx1X13TIKhbEIRE4X7bQsxRbesLY5MjSO78wNiyBI//o
ETWzHPe9lXcjOF9nacNBmP/y+1S4LFT3HvgpVyIdmzUBHvbvY54bu3Gl4mBD+jl+
RE4oWm9H+RAhiI6hG5oqMzNeJMqPo7c7Eh994gTJ5Y8kI8699slBDivCDSs2sG4T
Co96kKaGgEro7h2vCtFQ87Mz8VdR57qenIhYTKFo1VFlzDglVti8ES2SQPOW7N+z
xf1bBhrxMe0YWA9HtA3kJmNQ9OpFBTxTrpRb+dRAW3fCrjFIwo8I81DGarCokO15
QIMTrzO0NuVkk8L+5PuEgBZ8UVoEDAwII71bj3KcXwbXgs3nfPFrjQombvjKVmPI
C0O0dEzWK7xdI2PjGj+wt9kpSg/ZQhLK2YaZcFsoT/sQcorjchENhUjk+yT7eslo
yQ4HNoS3ubhHNGBzMn0DxomVUW0TDd0Vub2/IOC7QfNlA5E+CDlhrQldDlhziLMH
iOdP+Wm+3fpQQM/+iIF/+skNszb67Zit3/Ea4wB2VJ3YxqKFv/65n74cAOSqdvi3
3Btmw+ARhiLZ7jWMntVimfGGriQRzLGgyHXzOjS/PHZsOB2Lzhq8GZrJMOaZsH+T
pKfj7ERVTZy3PaReIqbyczr+sKgAcqH/upLkyQN0jZ3iO1yNPnKaol931oH9qHB1
CUO21ZlCa5Z93wKZ7Kuipgrk6yxtuCYj3/FW+Q/OhBWxtCNHCNMqbRAqm8zA1Zt9
ero6UOx1YCVyI0doNodNx1h2casLGHBxtS5BrTs6OxEED0suhnZka9mdU6PVxMYZ
h+M6AelcRMkCJ0+QEV6n5JQG8bSPAs4OkWJumRcW+YRy+XIH4gCMyNQ9yDdGQNSx
yLILsNyJsvajLs6HHeUqDMucffnWQJE1Vp79uOt60tHLrQr2A4CNgHXiql67eMbL
v98d1tgZrk2mT5Z040QRZskBuE1GxAfHwbDpE0LLkKBXIwJSo0U9Ka2JMrdKkv26
`pragma protect end_protected
