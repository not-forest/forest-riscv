four32bit_inst : four32bit PORT MAP (
		result	 => result_sig
	);
