clk_pll_inst : clk_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
