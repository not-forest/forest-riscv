-- jtag_debug_sys.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jtag_debug_sys is
	port (
		dbg_arg_bus_export  : out std_logic_vector(31 downto 0);                    --  dbg_arg_bus.export
		dbg_clk_clk         : in  std_logic                     := '0';             --      dbg_clk.clk
		dbg_cmd_bus_export  : out std_logic_vector(7 downto 0);                     --  dbg_cmd_bus.export
		dbg_data_bus_export : in  std_logic_vector(31 downto 0) := (others => '0'); -- dbg_data_bus.export
		dbg_reset_reset_n   : in  std_logic                     := '0'              --    dbg_reset.reset_n
	);
end entity jtag_debug_sys;

architecture rtl of jtag_debug_sys is
	component jtag_debug_sys_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component jtag_debug_sys_master_0;

	component jtag_debug_sys_pio_arg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component jtag_debug_sys_pio_arg;

	component jtag_debug_sys_pio_cmd is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component jtag_debug_sys_pio_cmd;

	component jtag_debug_sys_pio_data is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component jtag_debug_sys_pio_data;

	component jtag_debug_sys_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			master_0_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			pio_cmd_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_0_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_master_waitrequest                    : out std_logic;                                        -- waitrequest
			master_0_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_master_read                           : in  std_logic                     := 'X';             -- read
			master_0_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			master_0_master_write                          : in  std_logic                     := 'X';             -- write
			master_0_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_arg_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			pio_arg_s1_write                               : out std_logic;                                        -- write
			pio_arg_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_arg_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_arg_s1_chipselect                          : out std_logic;                                        -- chipselect
			pio_cmd_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			pio_cmd_s1_write                               : out std_logic;                                        -- write
			pio_cmd_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_cmd_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_cmd_s1_chipselect                          : out std_logic;                                        -- chipselect
			pio_data_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			pio_data_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component jtag_debug_sys_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal master_0_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	signal master_0_master_waitrequest                  : std_logic;                     -- mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	signal master_0_master_address                      : std_logic_vector(31 downto 0); -- master_0:master_address -> mm_interconnect_0:master_0_master_address
	signal master_0_master_read                         : std_logic;                     -- master_0:master_read -> mm_interconnect_0:master_0_master_read
	signal master_0_master_byteenable                   : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	signal master_0_master_readdatavalid                : std_logic;                     -- mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	signal master_0_master_write                        : std_logic;                     -- master_0:master_write -> mm_interconnect_0:master_0_master_write
	signal master_0_master_writedata                    : std_logic_vector(31 downto 0); -- master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	signal mm_interconnect_0_pio_cmd_s1_chipselect      : std_logic;                     -- mm_interconnect_0:pio_cmd_s1_chipselect -> pio_cmd:chipselect
	signal mm_interconnect_0_pio_cmd_s1_readdata        : std_logic_vector(31 downto 0); -- pio_cmd:readdata -> mm_interconnect_0:pio_cmd_s1_readdata
	signal mm_interconnect_0_pio_cmd_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_cmd_s1_address -> pio_cmd:address
	signal mm_interconnect_0_pio_cmd_s1_write           : std_logic;                     -- mm_interconnect_0:pio_cmd_s1_write -> mm_interconnect_0_pio_cmd_s1_write:in
	signal mm_interconnect_0_pio_cmd_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_cmd_s1_writedata -> pio_cmd:writedata
	signal mm_interconnect_0_pio_arg_s1_chipselect      : std_logic;                     -- mm_interconnect_0:pio_arg_s1_chipselect -> pio_arg:chipselect
	signal mm_interconnect_0_pio_arg_s1_readdata        : std_logic_vector(31 downto 0); -- pio_arg:readdata -> mm_interconnect_0:pio_arg_s1_readdata
	signal mm_interconnect_0_pio_arg_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_arg_s1_address -> pio_arg:address
	signal mm_interconnect_0_pio_arg_s1_write           : std_logic;                     -- mm_interconnect_0:pio_arg_s1_write -> mm_interconnect_0_pio_arg_s1_write:in
	signal mm_interconnect_0_pio_arg_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_arg_s1_writedata -> pio_arg:writedata
	signal mm_interconnect_0_pio_data_s1_readdata       : std_logic_vector(31 downto 0); -- pio_data:readdata -> mm_interconnect_0:pio_data_s1_readdata
	signal mm_interconnect_0_pio_data_s1_address        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_data_s1_address -> pio_data:address
	signal rst_controller_reset_out_reset               : std_logic;                     -- rst_controller:reset_out -> master_0:clk_reset_reset
	signal master_0_master_reset_reset                  : std_logic;                     -- master_0:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset           : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:pio_cmd_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal dbg_reset_reset_n_ports_inv                  : std_logic;                     -- dbg_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_pio_cmd_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_pio_cmd_s1_write:inv -> pio_cmd:write_n
	signal mm_interconnect_0_pio_arg_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_pio_arg_s1_write:inv -> pio_arg:write_n
	signal rst_controller_001_reset_out_reset_ports_inv : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [pio_arg:reset_n, pio_cmd:reset_n, pio_data:reset_n]

begin

	master_0 : component jtag_debug_sys_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => dbg_clk_clk,                    --          clk.clk
			clk_reset_reset      => rst_controller_reset_out_reset, --    clk_reset.reset
			master_address       => master_0_master_address,        --       master.address
			master_readdata      => master_0_master_readdata,       --             .readdata
			master_read          => master_0_master_read,           --             .read
			master_write         => master_0_master_write,          --             .write
			master_writedata     => master_0_master_writedata,      --             .writedata
			master_waitrequest   => master_0_master_waitrequest,    --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid,  --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,     --             .byteenable
			master_reset_reset   => master_0_master_reset_reset     -- master_reset.reset
		);

	pio_arg : component jtag_debug_sys_pio_arg
		port map (
			clk        => dbg_clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pio_arg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_arg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_arg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_arg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_arg_s1_readdata,        --                    .readdata
			out_port   => dbg_arg_bus_export                            -- external_connection.export
		);

	pio_cmd : component jtag_debug_sys_pio_cmd
		port map (
			clk        => dbg_clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pio_cmd_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_cmd_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_cmd_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_cmd_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_cmd_s1_readdata,        --                    .readdata
			out_port   => dbg_cmd_bus_export                            -- external_connection.export
		);

	pio_data : component jtag_debug_sys_pio_data
		port map (
			clk      => dbg_clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pio_data_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_pio_data_s1_readdata,       --                    .readdata
			in_port  => dbg_data_bus_export                           -- external_connection.export
		);

	mm_interconnect_0 : component jtag_debug_sys_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => dbg_clk_clk,                             --                                clk_0_clk.clk
			master_0_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,      -- master_0_clk_reset_reset_bridge_in_reset.reset
			pio_cmd_reset_reset_bridge_in_reset_reset      => rst_controller_001_reset_out_reset,      --      pio_cmd_reset_reset_bridge_in_reset.reset
			master_0_master_address                        => master_0_master_address,                 --                          master_0_master.address
			master_0_master_waitrequest                    => master_0_master_waitrequest,             --                                         .waitrequest
			master_0_master_byteenable                     => master_0_master_byteenable,              --                                         .byteenable
			master_0_master_read                           => master_0_master_read,                    --                                         .read
			master_0_master_readdata                       => master_0_master_readdata,                --                                         .readdata
			master_0_master_readdatavalid                  => master_0_master_readdatavalid,           --                                         .readdatavalid
			master_0_master_write                          => master_0_master_write,                   --                                         .write
			master_0_master_writedata                      => master_0_master_writedata,               --                                         .writedata
			pio_arg_s1_address                             => mm_interconnect_0_pio_arg_s1_address,    --                               pio_arg_s1.address
			pio_arg_s1_write                               => mm_interconnect_0_pio_arg_s1_write,      --                                         .write
			pio_arg_s1_readdata                            => mm_interconnect_0_pio_arg_s1_readdata,   --                                         .readdata
			pio_arg_s1_writedata                           => mm_interconnect_0_pio_arg_s1_writedata,  --                                         .writedata
			pio_arg_s1_chipselect                          => mm_interconnect_0_pio_arg_s1_chipselect, --                                         .chipselect
			pio_cmd_s1_address                             => mm_interconnect_0_pio_cmd_s1_address,    --                               pio_cmd_s1.address
			pio_cmd_s1_write                               => mm_interconnect_0_pio_cmd_s1_write,      --                                         .write
			pio_cmd_s1_readdata                            => mm_interconnect_0_pio_cmd_s1_readdata,   --                                         .readdata
			pio_cmd_s1_writedata                           => mm_interconnect_0_pio_cmd_s1_writedata,  --                                         .writedata
			pio_cmd_s1_chipselect                          => mm_interconnect_0_pio_cmd_s1_chipselect, --                                         .chipselect
			pio_data_s1_address                            => mm_interconnect_0_pio_data_s1_address,   --                              pio_data_s1.address
			pio_data_s1_readdata                           => mm_interconnect_0_pio_data_s1_readdata   --                                         .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => dbg_reset_reset_n_ports_inv,    -- reset_in0.reset
			reset_in1      => master_0_master_reset_reset,    -- reset_in1.reset
			clk            => open,                           --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => dbg_reset_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => master_0_master_reset_reset,        -- reset_in1.reset
			clk            => dbg_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	dbg_reset_reset_n_ports_inv <= not dbg_reset_reset_n;

	mm_interconnect_0_pio_cmd_s1_write_ports_inv <= not mm_interconnect_0_pio_cmd_s1_write;

	mm_interconnect_0_pio_arg_s1_write_ports_inv <= not mm_interconnect_0_pio_arg_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of jtag_debug_sys
