alu_srl_inst : alu_srl PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
