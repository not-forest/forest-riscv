`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dIqfQ88RLECogGhksSrpKy6/MytZUTR8o/yTO3jzPLXbOK2CekZ7WZr+n15kl4XU
Vrv3FgaxkvQADVTFwP1klv8VbgWWVK8i4AazJ/Kon5Wn+YG1wN/5vJ5gqyIB0ry4
TOUxL6Fn3riEFMaWVupGi271b/Bh7z8GxzPrNIzXg5Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
85/tnDiCm9/n+KvRVDYAEaD5hBqmD4io3oJ+Qv35sFOGaGI9MM8aOLV5NxnIF1t9
FQ7ugzkA91XjPCBLkyHUlHHWuz37OsJEi9ZTxaI+4eHrWU53vt5e6DyA6RyKev4m
F0azDVrZyuNBPtpAoeBU4TjNPy3Y5GQ4LavocP5M9wRS+AHlAOPBzc0MTuOGfiDU
Eak7jt4TBN8O+OibPFppjpcXndX4abi+d5JtmnWVM2A7gD+TYxgV5+/rIDj4ZRZ+
LD0jH0c46ft734KyU0+BKBZMUYJhowxVSi4/uL23UiFbB2Re/y7W/105kaan2ivJ
lzRD3NeGZ9kl/gqYkGZHge7/txBuQcxl5ZE5zVan3LMERwWlHMn30Cmt1djsnus7
0IwLRAVafksE0JIFXevQsg83bbLZ3QM6L5MZtLWGVyDNNdKic5N/y7c2oDOCQLoC
1/7U3KQzJ7ogKSiaE1hquDHY6Ism1lIJ04WBxkaiEevszJfHpw0s+CsN98udU4Qs
bY7dwfLV2bZOd8hS2s6IYH3QKM+vDl9IPV3fMfxpbLspezuRbsHKjwqOsTpNTf3z
92lwin6QPqaeoyCXowsB7SJkSHSY2kvVclmmWK3t4ToA8mLqeEnVW0+wu7/ebCIy
zeeknHglwITbqI10nY7eKn9uZfTtZeDTDdMHZhxzBNfYfZendXFaxIcx/l4to7c8
qRJaGeyJhBwqYBebmiogfifFVHfthcvMhebUJ8TdpUrJnRCXsHaK7WERup6HIdd1
716TiW+Nb5X12Xn9jC9WsBHHG4Lx2IDsp2oe3slouBhCOSmrhqDTVYLqiPuFVxX4
9VwU7Ur0OFAAmnsFT4JoE8UU3MaxQG69PuUBtJ6heGjfOlMBPDeSy6CLElf8NiF7
8Vq85DNkNmm57ZlIFacMnR3J8v7le1BQKtnydSVs1yEjhKjcZ4CR0DJc3DtlImLD
+hBUlTFlRePiG1rcEF9h+9cgK0RPh6l89+7zGisfHJ+om7nBDiGe731B4O1xEqm9
8uWvl+ImxxqQfOErtg8V1cSDT4WHCYlMqdBc8BwE2Id8J5JVEuOE3wdNavvImyK6
6YMmNuFTVHb8MF2MZ35ENHq7wUuJWVEq1CYadbhQRlyrw1Mel/899bqhVOP77qQV
C4wuJqdgeGLFJ1iC0lcYMAEA8+OBDWOq1/hA+qYvCO+fIZU8zESzgOP/vHU/7Hoh
9U31U5e/jYuVqE+VwDxp5LzrdhEZ9ocNmo1gMlc2LAuaRk+dDJ0GbnAPMMz0QPAh
d6NUtcd+5qqI2xrGkuLppZgiEmGGjOBthX3kZaIYG6MuBiZkS3DafEvtVuWtes48
ZFuNCcShvZwJYBoAHJ8w/vFqG+Sq+mRDiuLaGjvGVCQewTXr7s8LiWb2l8dL1Erp
ZesF60/fuds8rADGFPeaaUbpgrQ2hJO7BKsYH+dJl9Xd2AKoqDbqwWwqPLDBpGLv
oMeoL7R1f2X0CIYT+8Hc0cv8LbW/qsmAT8xE5jvSSlJ37vITbUmnpRHICZ7B7j+Z
tLxTe4Sm3TSqzilK7IZepJSH8n99YYP7ogez2oA0dtCKhmCdA8XLJQHivBzhwb/c
T6Xtt4cp3FVFUdRgIHSZxNxALCbnPnmgLzLUBGpHAgp7GDz1mv+FL61jRFUhk024
JbFmAphFJ6vmpKF1o+m+B+e772oBaL0tRsYetUSsmh+gU9oM71sHlIBBWAmwqql5
Z3YFLl2zC5izWY+6BdBtamViYkr8ctSglf4tOJCzgTj95mLsbk15UjmNT6rGKSRP
fLaiIvu3FcJsm/6MnBKFRYxgqtEwPgTHqGikArqQM5UoCCtEn3sJtrQrKqFndHcJ
QDi5kXgWa3Ix2ZEKp45ghCS6ri1zTiryC0AAX5hpwFPI5tSNPHF+6lzTkavlU8hN
GWSBvh1dM1iKDCo7brQiAfBC/2ebfu86KM3fuwrIR5n3YYpqcgygMe7iJHzsznWc
x6Xkc33UDb7Gl6u0QK4CIIQc/l/Ddgv8DUE7DtbIPyjsBMmRIvkPGyyg9U+y64U4
UzflHqH4oIFsxKK+nq8ZE7q7MVR6tRzvxz4pdrbtHIhIx1r4dD6lxTT7i0dJ/B1c
QELc4gnAIVH94zmhSGWWduL+Cy+2hQ9D0mBwBaypGGN/bnsr4v5UICs5vCUbCbnu
fC4N0UkVYjNVR25Y+rBJXc9iNpDqNtgrOt0T0gBuYTVlv9Wxvq2JTQRtvl0VUl06
2gu1yiWpLbde6KHRb/JAFh9FBJKF6KKMXFf5JEt+T4VJK4DW/dOt7+uD01W2Dt52
35i8KhdyVKdt2Y1YtFQO4OS7uapm3x2Mx97NQ7G73WL8IpGZBY7ML1XIb6XNDdMM
m5KvyBxpgatpefbA4Bds+r6gqHyw3bTzDlMqDWHYRGfJgzcyDLiUBIA7Lu4ntyeE
SM14YvmY+snKierHkmINH23+KdqQe/YABVCOFEIUC8CMa/C/Gr0N20C6CsSlXxfj
rKCmmZGpZvIoiu8oPS/s4YQSIwz1xQ4h8Ru2vz8l3dv0jtTDGo++S2/WtF0ELmR6
wBIW6HN2lFVGGf5iT+VQsBMiybWTop4WByUTPsnPROvEMEttDI61KL02N7lDMaXQ
eIbmkoVgRCCvQh+Gst9fYnFny411yqgYwmlrFKDRPhNSQhummk9CFgzMYAdNPyzf
Z+JJOvTPqTG99IuNRZVxR7GymRZQUZhasvk8/jwrZhZPkSzi7ss/UlA0SW1ApNI6
/u97w0dMFTM8m75tV85YBEs5tAcnazpLDS6bo8W88On7L72cDLEZZH7SCblmSl3J
yGE/JSj9CNGf7HHFXu8l/LJEjAuKhM9+rI8/zj2I2lrE56fnm3+k/ixoWgUfra0f
yp2SVa0R4+k6RzT8DSj/yKLKOKaQhkEcxqW41Fk2kWTR68KV1nljoGYuMEqWpZe9
DppPkDHDfSEXq5rIx7ihIHeVraJQaf5k4xu2IvtNnH5GfR8cd6FaIro9GfU+awQm
jGwmc/hhJTKQb9hfwAt9p6lDnGLG0d6KiwBRBZuoAbakQRxcPu64Ukd1N+wfyowv
SdQnmjLst2NkvQmGFnKFHdDrSTeILcbPEj+jusBfKVfcRYgp/9H77zNSCW+CaWzJ
M3t9lWor3UqQ5NuRF3TNodc3/M4RoNrSMgECS9dTd9zmcxaIthvY3O7R4j6UUoFJ
QlymDF6ObYn98IYr7JjtBAOxfWlP81SEHN2GAfBrosutnU08P/DXCurahFvxI+fj
902XEtjZu4HYsgC+kIew444uqMzPxBjkLN6vzIHhqlkH/xf0aEmzyY46bRCC1k3F
l3zjMmGbMrqQC4BdL2BvhR4DjwwKHG0Gfpzx/8hgsbJ56XYlw2r+DVMQCWoC5V/q
FJzOMzolwQw4lehIp18efl8yNouNxIGQbMXuQZuhl4ikNYHKNf/P3zYTtwcwAv89
LLTDG1QM7CnXUEzvZh60HTtnNgt9XW6nRD29ZkJ3rVhx12CadMFBlYF7V1Q1fKci
Cr6AKJsR/XxgAusyzSVjMB8j1P4TvyXNmW4BMXBsnRVjTRo7VYTcZq32b0+Lyo+t
qzv/jT1rPlI7x9dUxpgQjXTlxHLE42kpiRcT8DIVqQYhFhazCN5Qx4DtzLK+XsfD
hTDp1judGFgZpwjW1Hyrks+xafNFdwwU2VdXt1rtnBo9eCTTbW8bnVWK9wFIJpxP
uJ2SKntT26IgtcAd/jMBntrrUgQVRA7lL5HkeDH6PXFXByR92nRwDiBCpNLBo2W9
GP0pKA8mUWblVQOTB/ODODucasHsbHM3AH22TlnnV6WBVGEeTM305oZRiMgBh4Tw
spUZgi9H/JeO7yf61dBpODzUdi8dX0x5K8omBdonesb6BD5xINken3qHhWECdbqr
5lSfhd3SQ2aMy0BsQ67yoRMMefytpUrOhHuJPMzwGqZK1R4+EpP5HSSaeZ/EfLIO
2Q9aPOtIauBH7v4X6TgExpaSzSV6Ds2HTL/Z+Lnz8TcxXVc7nLcUHrMvKfRfi/5L
uNRgOFEERKdFkqjBwQ2sUCdNoSBmdP6uSLmI22c1zG05fq/D4hO0ia+NePqiwS4G
4UgQgwnL/JU/7t1f1D6VyEsEbbC8yn/q+1axeC1WH6DawNMth6xfKncImsZIQxDv
P3u4GHbD+BNqe51O1WHwmAZ/TJYBLj3Nw9sW15Q0MXKZem625xF4YiR5X9ryzjA3
tivUhKoy5fdD1i1YZUceXHBRs/nBoWZvvpo55FD3zRVVca2wqpH6KLZCWlqyFowp
ony5rA/Cr0WfFGROHtSo+ijNyYosenFq+X+LYVwII1/uutXIwAYR/YAa2pzMw9Rb
7qHfEEV2qFk5G5nwXv5/niPadZDTTAFSJ25TUP6Nk3OeQ7RJnKLXIJLaRZPs7xyR
LK6KDkw2maAOIyQiyQiFJPOIv65/kKYEKnqJ/NkBLlDFTh32p2bK7orQN5VwsGwr
TNdr++G8CGOFC2T4eg5uAOvHX/gP8rMZiW79k+assseVXCHcsrNclwfk34xnoqYH
cY2Nw8LDw7Kr/XAmaAwjwB7skEhfp3V4Su+A/an7ig04B0PxPdVNDzq3Ucvozqet
mB1D6Xpyt+iEngm4kZAwQEoW706n0LOHlGnddgIxgSFBomWwO1sVe/xLTcVVE2gj
crNldRXsPiEht4vfkgxdxEYHMVaMFP4kNKbzBbOUGQy9SHg6m2DVt6ryHkvK5yEK
Daxw/XlydP+qvg+6kf+m3hhROHtVCVgyH7wigBaGIzvIeORw4wVDup6PJ+AB2KE4
jSoSNHYawKWZjhEV/wu6t0VIBjIpEZw4AXgERO5DN3cR67Dq9QTOTrl/rwjBS1px
7Z/3Ziij0W1BWOVhSjxsOLwyNGxj4pGYdVclVdF7ueGtXAIZrg53Rd6Eve0d7lQp
NUXgKx54JKytNcXTY3JRAfGduEEkWa4x8up/2cXYWLEut33qohIrlvVHWu03GBjT
1FX+HsqbflJHc4dchMhEMZnmDOnZORAT2qX4YfB9FKbBuvqM0k6zuDC/nwH3Tg8P
pNHppA5ZKJqF2/VURXcw0IiuhWHzgCLFXrMV11z6roBuAb/rbkVv9puqQVZ7KghU
WUreXU4cuKvlbdE3jcyDdIiwBjDPWXbkJ0JmYDnl4PhUvCDkLmi9qTyt38VrTMy5
UHiXk0oGiMKxky2ieh37/Dq6cGGev+d/bIZI8iALZSlP788BqbuoVHWUeevmbfbm
YK9KceTtX++aA8Le/ASTjEw24QtEYSJC5EXbDPolHrbil5D2WYA0lAMejMWZQij3
TYfF0X3FJk/hOKFka+EUWcKTuKLZ+fvhfNE2izgaDslubOWFJBaV19qrHefOdARu
FOcsNGORbDZRzMfGjtTJAhLfwj86Npy+KNbnw0SowLDeKV7ogQfIafNMQmZsPVf3
oMaIjXfZy36PAIqIV9Ooi/DlHshGEpozBD3ASkgJIE88ugWQkdrWIbnuRzomXrMR
eRrt4SOwqgd7Rs+JJbBz+VPA8G1giylbb509uRZKGFSYjY3OVVmsammlbC5bILO4
RVnZxADZQzO7i10SPUrWkrFfMmrYGgIR+GVsnh9z5d5Vdi55prQmYPLakpcPW4a3
xXrfNaSshEC1DrbCJ70KvhYoOj0ivcyM/Vv9JVQftPYqHsr2jfxRFo0+MQIxnpU9
LcCKigzCrJdZnXf2CyBqPfT9NKT0u43WeC27jDAk8Q0g3vnfzMehpftl2YVeQSaQ
Cvp9xIR5jVfQ/cJUSyIgGDNjnqP7Ligs2++68Rd6FVni6vxM7/wwhYYHbGr7D9LH
cEdMbB9JOn01TdQoXvRLBJKxcZtF3gsz09yoecDbwAypI81e6o26OEgeEOvIb7cB
kQl7pUwkxqXH3Fi27nsqwf7ykWHq2wQlk0BaxaOwZn1jF/I849Hi0F34Oo6xgcVP
G6kZUNjZXkd2rXG2IgNsE6qOdFaDFzd/KKCzL18qyW1tZVsUrtJBZui173UN3YwM
2O/cFjRlzy+elNkIWRRXARE938eugOGFEkszenLsKKwEWxrQRcnGEkIOEFNhljyl
a/Lku4hiYcyFkN7tGQnl2Ko7+yx2MBCsY1EE14jD08pnnmd0qHf6R2UGlLabnx0c
8qxr6oiPvQ7hGKueR50h6QpU71Sn9pk346CrK9i7i82PW6T+N0FhXcDaDJPyiV0b
7SPI/8Rus6i095jssqRqwye4MQw5cUt+uI/ky7IFDyK8KCOnF9WJEmzx8QPIROgv
OdoK1VpCvxwh0lgR5neDbnkxi1101LsW1y4sPjlkJflKJg+zAsXUaL+ZMttjmf6/
D2tVUDOeJZlxWVdU27rGfbr2dAXz/mDPY3iTtoXW1zD3w5S4iwrnAswmUMJT3gG/
cAQ6br1FdZVax5p7HuoDU8m7QyYnbbni62YcTSBb2/Dc6UaUmNWVmg4jkLI0bTQ2
TsqpgZ7ISLTFwNGvdNDUw8fKhoii58PaARG+Y8P0Z1BI+BL7wjv0TmFYj4AMeQX0
VBpZ1QJM6cwAqttjEh/uq5/PwfdoNfKAXnVejGX8jw+TW/WcoXjw4BCr3Ydzz+In
KRL+MZZ9Az6ZcZkOnhegrqJCF0CvO/Z4KMGbaB+3HPuM7RGCcxS7DN3zpd/B3HjY
QXdhQHaw11Q+h/YLij6t1i/oivrs3MyLTbl0Mmu2OYSCX4InNIsEvTaRZrAxRYNH
EIxYp39vo0dnL7PNNx/YLlxh4MZJmxqwbSDoLg0a9BXTWD1NIuA8O39lzZ9kG0rb
XJiXfzjjOGRU98IzvlaBLyZSRwDVkG6OGbOzLxOCTPvrCxZUYjm2KMsgmovVOFCT
FUEdccLj4qrt03kR1J81Ccp1qijTectj1BjIpDUjHpAVYFuSwXBfGtIla9ly+wwZ
sjZ11yQXWJFf7D0/lrL0lHLXvq04ZSmZj+f/o3KJWog4icT0LN+1fdspchd+ANUe
RUONgLojwzGwbtIlTszMOn1bGdp0ADjD/WcUJWPhTyKgqzAbSYP9sUs0H0hS3zoh
4zjWwcI0K7WUa0+H4Qg3RPZPw6GNdEWIDu8ns5fso3awtGaJKIDGSuqLzksYalZD
KlVHhCRqmh95EEXawQVw45eoQR8NRA4gO/hJbSJHJ9OcCgEJ5Bnj9mnfu+3qgdV3
lSLj4xak7ssS33LowZpkeBgmt94PN/pZlPIV3pWu6zQj2oQ5cJeTCfObg/7cC5qy
eD4kt5PMHKWqzzsK0QyUBRIYCrdKbshoC06SQ+s9Uh0ynRat9iytjSoqTPM3UsJU
bhuWQtIHRJO9ICwaPwU1Cv1fU2NJli8mOztPaIyn5DkT+SleJOTYHpoJ+6IRIaiP
PMwHPAY8mb0DfQlQn+9RYlbODe74y8x169yl7K+2yTVPI2PvMcC+GyEO6SL7nehI
Ykmf16nNkaYsoshPwaQkZsZf6x2kF+Cx7RJw4Unm3vaW8Zp97fOr5P9VK37oU9hI
R5i1pdSODKHTPGGpHTAyY4ueZzRLgffwcmrm55AQJ1KlEhm/wf9VLYOz80se83ej
YYh+Yd/mKJaDjn1IwDM1o3+mg/bTQMsSu59IdH/01zyqHcAOiiV/11MJOPd/Ki+S
X7W56Og9d4BXpkWbe0qWKRli0lZC5fseE5YG8ELkIuG6eyhE1XLJwawcoFlETk6p
rbEx1CHZuIGlU/Xew2ERIm8VzRX3fYMAlbpW59pk1/0UNEyD/q+nqSwwGDTk5HYF
yaZanfWTBCCgJtwQ4kUdjZDCTYyNf1p1xIkRGnd/wn3dze/+LdU8LMo0y4EZ6N16
dtMhacb61Z5HDHwwnpWx6Lv6xQoHBdI0q60sXYEgxlSAQhxdYCvEb5a7e5vOSBhd
XQvqmAGh0zM2A9g+yhYLawzNljpkwiq4brWFzGHd1qi0oUGhX85oUKECgMHytvFK
fCOpkzB53R3vt6+vIfbJACz0mZSfCw5Wd5NpQ7iPx1VBhBkSW0r27jsshtRZ5WPl
3BhounaS3UZGTjNklr9T/nLPeipWLe95B3wiE+7WV+IOaF8AKRoQP0/nHjEE7mfr
6HwQuMpcOskI+Q07Gfkr79wbaMgvqN1137yI9QMAVnfJmYnJivw3iy04uzbRMzyn
1gDxljh9yILjwJAa0bG4TWJHdO4WbgOhW3jkIl5cWugijbgPLfYXw8oTPNXbQmiO
7ctP5yMjxC1PGfUQWURtP7w76GYEs3n3mbCH05Udk0qBHj9sMUKu0wIEXnK+Y3hC
/l2j7higtzTvHtx+d3TeMgfT78BVEEmtVjs9w56lGIJEM+sxY62W/0mi8vC59lj0
ld6tISfgykIS8EIi8xx3duSoD7TQok+hWhSsASJoKKGMqx9mcXQuhgBm7wnPs1Xt
hRG2rn/yCUimhNsEblnkhhfPYjBeCNRzXO/8b0sn9sUm2MLeGYHZWOQlhcxuUH1Z
BDi5EJttl/TuQN8qkAttSDPXJVPjxpbtr3xbP4KKYWEubsOnbOyBKwGj8vW7NuUp
xhMRPzUvLccduedz/Rb3JBqfVV/4GhaU5RrNwru5po6/GgfENDP2IO9XJsmstanh
QVIlvtvA4YWNWmykUopNYkdxhzLD0uTjRHa/9GbrFMM+e6L1Ih87HbKKYZSf6Vvf
Y9ndTxCx5dC99qRcy9WPkjdrNojBk2zSEkOQp1ZxfT8DrbY1W5SWl993THqlGn8N
5q2zjzR/tPseUF6dBPm2LHHyXyoFBDnTrabGDYPiQRr8vYjtoysaxFTd3KZGIZtf
C4KWDKl2z6MPA8il17qkFCqZ3gVo8hgA3QT2C4o6fCgjiyXog01FsM72q9FW7cp4
/pmy/SxAeChC9TNUdHkTv069ZfrUf4kbnrY9SBwJrseYZaTJ8z/tVbG2jLpPHUrq
yvzP7VqPlSqZifq7trlAMW/FxXdYUHereoOr1WJZHVCoWuoKqxnsXngWvqajBpsN
tZfnDN0qZn8nFxIjZu7HBgGVaCPnNolQilCojDuQUq0tMyXU6Pi2RYNCkFq9RykV
UWrjt2+QCdTk/l+lVpMqHpC9tNOE969T9VKgZTGkS8oCIO7pGQbeVICZtSpw3JfO
pOMl1W3JssrP+hSUZCebkjKoqnvWoobt1e6QFnuvT+qzeyXhNuWek9o3OUE2Bzde
uQUUD+VATFPd6zTfJDTS1E9UcOe6XIRPwTSDBUqMBrupAzPjWhmOBxjCFDDU3N2V
AWS9hAhnKJc6sMTVuO14rt0nc+p6yxq6+Vr5i53MFfq+LYBegCcI2VLbchZsKtqg
01XpmSi0kMT8gAxcBVraGnUvgKEjzAFfhy5zNlvvIWDixIoGA44KC0mIWWwlUdDs
1KBy20gQO3c5gew9HFdJqKEzyxJlqBShnzYxFszyyYboShRyiyR1Od4KdFa85q53
WzpUaiXpWzxmsX8Uq30DDIH7JfEfJ+Bree5gGNLBBH+nBnl4/TFiQpmJ1DBA9zW7
`pragma protect end_protected
