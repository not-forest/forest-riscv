alu_cmp_inst : alu_cmp PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		ageb	 => ageb_sig,
		alb	 => alb_sig
	);
