zero32bit_inst : zero32bit PORT MAP (
		result	 => result_sig
	);
