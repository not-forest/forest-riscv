one32bit_inst : one32bit PORT MAP (
		result	 => result_sig
	);
