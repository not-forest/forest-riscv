-- ============================================================
-- File Name: pri_encoder.vhd
-- Desc: 3-bit priority encoder for choosing the source input.
-- ============================================================
-- MIT License
-- 
-- Copyright (c) 2024, notforest
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal in the Software without restriction, 
-- including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell 
-- copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following 
-- conditions:
--
-- The above copyright notice and this permission notice shall be included in all copies or substantial portions of the 
-- Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE 
-- WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS 
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR 
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

library ieee;
use ieee.std_logic_1164.all;

entity pri_encoder is
port(
		din0 	: 	in std_logic;
		din1	:	in std_logic;
		din2  :   in std_logic;
		dout	:   out std_logic_vector(1 downto 0)
 	 );
end pri_encoder;

architecture Behavioral of pri_encoder is
begin
    encoder : process(din0,din1,din2) is
    begin
        if    ((din2='0') and (din1='0')) then
            dout <= "00";
        elsif ((din2='0') and (din1='1')) then
            dout <= "01";
        elsif (din2='1') then
            dout <= "10";
        end if;
    end process encoder;
end Behavioral;
