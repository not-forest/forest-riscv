`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OFHhV1JdwPkm+2zt++q6rMSKsvR38sGLMKwygazbMTaelVE/FurdX4tOQ+15i6Ry
mHjgKAjfLnGER0KIVEEibdZZWM40U9U/+Z/+9t5Q6ptZkK9xsROj3wt94xFUapIr
UM1UR/hWo33tv6ZrYimrI23PApNAPi6srzHgweqSuuw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2848)
9vMxwGFk0H3ISkuTpvKAX1zhCuYAJUGtgYaUHRP7hwFDUBabY82XpyAF0cviTLjC
IKJHniLm9p/X1swD5DWf6RjsDwfYdVqDELA3thjvWPfDGtSiLiJAMI94/XDjLSLv
J4MDIxWeqXDJfteSN+cLan+aW+RJkMbg37eI2laPLEeWGlYOYnM7CUwNb1JNCXZZ
kUuc5PG34yxx+Vep0QfVLcLbj0IPNDJoZgWyEyyjsFtAEDFveqd/whoXYp/HAQ7j
WzcPFwHMm3dlz0OJKPRnA2Gi1oD2hX+C4M2xGeqhmnegrGMBt5Ca6sxRW0SSkIDq
APl8VjJ2CuhApyOL7pcqSjbqj5OvF2tx8MRuFByJg9NB3lqIFKrURU1seA8pBMtv
FtrRqv0lOvwKCjY3rRCt1XzPyMxT1A91Vahm1BIAeap7bYNMR7UtoRxWDYMt4AXE
k0mUA0GCsZDIHT64m6GJ7webqbatRzV50WCp5jpYU3sE3ACPkQZUZs5r31dfMg86
lMOfQmpJq3x/jn1GlTJGtF14LPpzCI9cL0YSlepCS6wnF8XS5PjZlWjmdoN3LQqD
yZ2ODPw5SRFbdwjITnwidVBUWet/fy/4ikNRbLn/AXjSDDE+oJOYV6sJ/NR1LggR
yARuZfb6pPuWIRLNQ65ux/ADZi/oDgd+k4Td+gITv/s1u4KiDEhrH6zFLAHcgUHQ
KqBJU3B5uXX5x6yrUziJUYs45C5lQ4EpWjj0RFlBy9bdexRmMJqyTc99TsXXSXhZ
/h+mhUe0j7S6i4Dle1hCVVPKhFLOMH9iZ8o9eMlFc8p57q5daPL1PbwdZ5qXwLCj
yNZvmGXv951VTNrnxiQlCqGa8DUhvII5zggm/hiSXqeYanAl2RKu5KZ8uGNJVCoG
z5ckkWt9T1GGtHAa+xHyNTUQaufY3Y6+boCBNiZtkBtVKK3ZGC+UmJQunfZv6QNs
Tc52bgHzwIT9vxyTNiM/qoosBuIHzfGa0zGdX99aYOIBtoxM1JvqDCt9FGUBSc5C
phjjRl33XAASF6s7D/HDpLhMRqaUFqqH3NmVQlmGLlW1NjSm1QUj5DxIn5kzRiLs
KwuPT83RlFB4L8JQqfz6nsuHbOCzDO5JfeSvHhb1YwrNZVXfzmauAAqSO51xWTKs
l1ect3Y8iIJEuEOj5soLSX5feQu7e+XpKos4zT+RMkL7ZTpkQNh7lO2i4ayW2Z9j
szuvSbavbD/V4Mqp8uc+bLOuVqWjdmpmlJ3J1Dd7+fsIeRC4FlMd2xcxaT9xkwWr
cRuKGc3J51u0B6xVB1JMQJ+lvTwhWabZu94H15EF5GMKzoe+oEXrxV+XxEI8Ts87
xRq+8eBv7jkL6lyWfVfrDEZfaBmRcatD4qDFGnrVpkNmpXlE+ygEry/P/hreDDb3
dVrRu8w9VR0WncU/UVnP1LsHQGQctQlO54xNLxrVtXYRhNoewXfThmgUbqKuE/nq
UPyqwpEkQ3qxyeTIt+SX998kpjKy0gAceNDXlkxK6c+z3LYkKuNvO/gvfM0Njecw
tg0+QHdft5DwltyfOlN2wk2esUZwH4X1gUOXYGu0rehRwGLvzHbAjfobjPtLvyNM
PFotd61tmn6r7qIVROG6rS3PbR4WbKz+d5zv38jFHQ6oJh5GAOFZuAWwBKKchd2b
hmne1z2aKbNMynG/4D1ESuIbRUiix8KarHHyGOv27IvMSyEV57kHg6niqWz5s2FI
Rs8QgqiVkCmd/XeRnqLKNBNe/jTNDoQNZGcYcgchfCCl37w8d2RjHq1IILttjFoB
z3aq4tOze7mB6r4qs6L9ni8p66bp5rM7zXmqf66lncVtjyGaxQ9E+B0Mmxnvtjth
m1NWjtpXneqQksMs2wgKdU6/aoG5SLi92a/PnIJS6+PozYK96vMDkA5SIjb3n6ha
zuLgFfBHhHJKSMtAZCFeS8OB+v9vQ/7lXLaQsON5H9ykor0M+TIzshlTH5YAnyOi
CTpcuyR9hYaBIRSJQTcpcDkm5ztSCqyi61NMMcS2krDQhCs487ycfgukJAyGpkr9
bAHPmddkvouMhb1PTBK7ysZjdDg/i308ZrdBTpca6TtMydkFifEcxRbDmcj1Q1pI
RSvi67Dk7ZbcylZxMvyUjH5Bl788JI3OITnLrqBKQEtaxzyODWPdK8caeJsIedae
QsLoizYMraCwTsgko6SqfsRnwwdUceiUEey4LOSeBDu9C5SFyntlCFvIVErf16Ds
15f7XnnLbDMjq5egQrzo/QI+DnSuIx0Pv4wpjO8ft4FTRqxiyILdChzW0rKblnHN
ElT4MLOO4iRENOBVnOAYwooEEtK795FNmgyrwIipYuO4Dsgmuw4B0Msp9WuUrr3y
gxE7OL4xmT1V6akf3C2bfL8qnSUXT3GothBb1AfMI8Hfl1S4cfdfoKI52lK23TL2
BEALX5Sbqlih7fRhte2Yjwc3+DYrnuFtFNFNBYnzDPrEtiBl4EgIQjsROBtihEM5
i3tCQTnYJgbNFaf7aG9H0m8ovvzVCDkI7N8O2sO1E5peqVvWqBfa+5LQ0/Aie8Qz
mUWilSPcy9G5yB3MAaHKH7PQo7jhrxsWH5zWgAuU7WDalUXo+Gpj8jnMm+IAl+B0
n4jANEMFnL7/pK/bkWxW3Z2yHiQoWtpgalgjG8q0VVLFhQqXrf975xmaU42u1a3O
rbO92W5Cyc5hB6Wr012m7XFhrpxrEhL/OymrEHJ5GY7MAFCSr8IyoABqvaRRhOOU
l1EouQuQyg+gNYtz8Ijl9UM/PN1mvPfdiqEg15cUtL+NQGyOrLxxSwSGhJ/uHnOl
CvduVyUF6eoBXZ0JVVVjhevI9UMlYOj15sHMXJ+q7Jp9QCBuZJdpvFz8rCi31BO/
pfpZMdmuM479DxI6/hfHyBW+KrqFFRKIXhs2bPD0Q/UYNBDh0GrkXJAhLIvejQMI
G/SKjx1xqiupBAB+Zo0XbF4wJ6rRwzMkHQ6wj30TIFVqrLpb2lQXJCmUPdKWjm7S
rrl20GjU+Gcm5aS8FNQkK2ypIcJUu8fBdZ9eKKOHv506d/USqJLxzZzr1tEaaH9C
XJlB2pMD+cY197sfF84TbJv90Dml+8zhvVQ/v2SSpNoC0aoeEawn3rGO1JObayXu
uCsCrkmYvP2Ox2idvfw8YjSxFG44NONHQ9BXJ365M5TDnJo6W9cH/Am2pxqQ9okC
Rk4D4Y+3YLLeNqBhqDudpE3+ms6gXNoBkhMwrnNfu8YvQrmdZAyzSps0ImAgAEyL
6B7YGOP3zFBzRKCvRihJCxXyD7olsUkfU2w7WeYYAY9JVG0X5ULwemMTZUIFhGm/
lRJgck6bKAQubJ5OO3YuL/wUSVIeN4AMiojUCjPp9dIJJk2YByhundAvDKl7e9KE
2cb4rsPO+HpMQmq5SMHG4nTGr9vNIm0rvULW6zHUkKgpHj7oGz/jcIIDR44bUpHh
rqK1jDfk/lwlCKdAe+IX9MG6N85o4+1JVM2y7iQFgc9C9n26H8CSM43SCQU7oHpk
g+bO5yS9HJr76ECna+iK0zMkCl3JH4eiL3F0hHBfvoU8oKOyZ7twhOoiTlY4xZ4s
lJLUKI2lCMfcWNXboiBDA4ovnQMdn4lvuIGdQNsorzNqyI39W46HEc1tGBMuzAiZ
keumPs9x+QPaZmZxDwo+hD+sZcxzglDag5++Hwe1U+d8afkrCSWkMa571GtxqglA
L1oAJ2clTa14jeyfVFz4Ta7TP60l77fOd5ESeSXDBKhRSv0usOfrfT9QlLpel0ym
0GNKEVChhvHcDA57NDbIGw==
`pragma protect end_protected
