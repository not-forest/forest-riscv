alu_cmp_unsigned_inst : alu_cmp_unsigned PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aeb	 => aeb_sig,
		ageb	 => ageb_sig,
		alb	 => alb_sig
	);
