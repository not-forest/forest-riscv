`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KROuJi3tV5yByG7yWp/kCRoszkoJLP53gs1kmz+d4RlEpuQ0vDK+NidRSRE1Ampp
2HCFy36RkIRuI9lwcUX2QXYdxrsLJxWi+d2X08bAh0N/dm3k2WguouCvV9LhjLe7
dA1NRejKiE+he95Ftbo+LbZa8vLSfE1RNsSh1EXDpVw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 82944)
2Lwb0Cm2ZaUvue0UEpaBpKir/PSAu8x+fmIdQdvkzSt94Urc89trgp9ZFt7L0nx7
i3smCBg90DAe789yXw8zmKioy4kLNmGMREovbH7q5yGa1EHu/vFkuq9RLYCK0WYd
+jy0Jn76RZ8tm32++RDMouIWQgcybuJ9icSfxuvY0JIU5mXZPNdBfHqtLvBB6z/V
NSuu3gXZnl2lSVPXgKqw08xOacr+3qoFYGRNJAWWO1zUlzucVFKvFT2a6p0yuKMZ
zt5RCjFSiF/UN/YMkIFIbpW10KpxxnR0DS0wxx43CPPtkRQZr3tv+eyFpGq4mKzv
okVZKIRnyMl0KztlSrA8bi0AIVvFt+u/nGrf/1gAJVU8BD2a/Tds9l9Af/ey93r0
bb4OXirHZPl33/5lQBMySZzNhytakr622MfTE8xHxBggc5BjITNX69DuzcQDoDfo
N2raDcsHxOs0iCR9fASsD8Ui+FSoNWK+4lNyf/BrmbE+y6L9p3UQLMzOxbLjHu+L
FyKI5nfcWER73ujn4yBE/VMtBXZDmw8BFKbVA1UpCZxWMt7ozyyi3uPSSE9VfROy
LPyzyQouRueKt1ZNSLoTr0DtbP2mywudQFSfIMGW0rx02GlQykaZ20b6bydNVk9a
hw4KDuYRX9WUeV4st/3D8oAXjc51YwmihgvcNRdBwvDaLb3E0rQ8a/4A726LujY/
Ork44XNN9akZcJ/38q2v2kUhEhSjlg+uX2Hqry/O5Q6NQo77rI827kqVkIY2VHPE
6/kZwecDOcZlA0L/wejiRMNGyc1pokakjmd+CA3lZ2Xag5FMPjFJh570wLLf+VAG
TWHFTuJMrXQYrLUhu3D3yKEPufwpOYGIYaGUcACrQndWn+ddiEA1fU7+QSkx+3Ev
UNKkXlbraSac9ZtTLhBQnZCHEAiu0D3aAoNKX0cdkKbGLq+ypHKHOmN+mN7eiSso
shXH6dTjQ7bl8yN3yhLv8I2DlV8+PHun8vUO7EThlnbLS1yPd7bgr8D1oG6Dmus4
AK7btuIskrGWWJ9Qb9e26O798BbkPN3FATn84oXL+emRYKrIxCuKmKkWtujVZBTL
6xFxtHSpM5c/O8vesmJizSCYn78kVJCv/wQ1MEWMRqVqQz2nlY0SuRdDwYP7iJKN
zGdtbh4KGsAREBp0zt7Ou9fiyTBLHR26i4swwHwLqUH+rFzctlxXoNR4EttHSQoa
jU9A+bSPe4l1cALcsiTjMBW+Qhpuvft0hfdHnkILXcuI7sehZ1nwL6eSYzn4PJMO
o4aMkEaOLgZiX3hre/kUv3phlgpgJRRoGeFUqsSEOm/cTvGFTHwOD9nvpDVxSYlv
9zow+dwyFFdPhooOShI4ronXARrB6yasAGjIMsEDi0Qr/ufvjVVKBTXnEzA41OAq
Pr8FyDFZHg4ChWUHll04KsZS5TcRDTY7GPn6GqOy5IW1/RyGDq1HdgJGhSIU7I7s
zQNUlwkwN0/Q2M9RrF7bnJr+FneC2UDa8LYnBnS8VKowMV4I4qyLX6c9vjzhyA59
DrNkQYH6nc3OCbYYOvbOkaKJXGOEaXEDW+8NnOlnDDSBydCrd0Ck5GVJCCGR2kF5
pp1gX4TrXl1jn45vxP1PYgP2DLlncqwFIypdqExSCZxcW7YbmTSYpMSyt7MbpQLx
xcF/BmM/1kEiOG9mpBYLCXyxRtaCHbT4pdmYOw1sJUlDG1VXxcoA2E+uWfHGN+mV
Zgp3gdBnHRubum/UecrfqoO8enHgFMFNy65rvzmXVfGz1nJMw+iRjmq6FgZKcYCw
3TJYhl5gUbP2ixJuILiYV89aNWv9RzeKydKvIocURIZ9D4d9ncbqLrs/l1PZRMl+
PbbODRmSMlItOdBvCSCvHp7w98BcRDcI3fI7zYy9tVkM2+8wtchhHe9qFvpR6ufN
oFNRFNNqchqTyhr/YH4b/FiCeh1KNTYFIt/ob98kv/aeVSwBIN4QYUymcdFav4Mu
sOQWWXzY06hrQRRboGaFTQ0Sf/OuQb46U1meCcGdSu+GvS525TVZiV49iQm9t6Lu
e3QVrAkOB2eKucs6+Cmh7piALJo9cBdMnPKC41+O/+G4SiIiEdqFUt+np6kyyLWb
ZZuzyJrKMp2g8ConfaTkMcir0g47hrkMYGR49NRZKtkTD21knw16LWOUQ6zceMNU
lJA6bpUZDXnLpjZCmfHWclW0IUDe4FwbuqqKUHmUzadGJ9Mg2JQa2bOPAmEuSo1r
ZZswDZqDj3A5jwF/UACxKovJxUgRUk9SPhDPEqfgAsnwsp9Akd3ckW1FwzigOvT8
6FV5GjrhYcS4k8sCSRQft13Rudu3kxCbEWLAZfSALCbIkJopFu8PnQtWHkjVPRd0
qNsJCohVeEbo+bkPVRPOh8pqK14oB1XsDPC6PoGeSqUn03AC03R7IsGgvyzF2a2n
ZzDkzaFGZgZ72EJd5rvgxrPwfe1oY9oIS10+NtpzZHO+eLJNOvE8NTtY3QFZB4OI
XXQAYboZvVQnlkoZr/xGKsswU1vrJ8FiYEiLrrUqEvF9L6sU+AuyikWGy+RKQLSw
eJ3eeWyD7s8TQSrq18BVKgOldWwTIDO2mPRV0wrWl10xdXlPWxUfyR0sqX7z85NH
3rJgyRmtn4AbT3lFvHg9loWzoso+Wpw3AwwGUKMQXRWt3oim7f+BNuvUGB9oryw0
dTHUss2HSnYinWtchCG/HHP6kHqz09tvvOwpQq5OkquI8H8rvk1eu+PvyeLkFhSd
b4rCdm5GLu3E8VTWlHWJNHRMVBxP8kOAnJJiz+K68wTCtRzBBmfsSHidf5tOptqC
SxChuYcXoiDh06jCm6BUFBmIG8u0o0oKVluocFUHGoTgO3dwld3j4CU/AEYk/i7R
G1vXfznUOALSWyp7twH9AlZsS1RCM7CVp/cdTcvy+nyjitC2v+RyWZzVpTW/M5h2
RW5fWPnVcjAE0xlyY/xiFosT6rbuwsZCV5fkK0KpziQJJA+lqRUF0x/L6auoC01i
xy7SmZyS8yAtxwtdSgefpH2t0oAnVPYUs0KCM7e+XBZdoTaSX14kca9dPHgQiN41
geh6e7fajGDywo+BJObHWeSbGMBYVn4uUKWlZOTVQ7SW/efKvCUYpHEz7OVssDrU
hXPhRyUm8JhraJS/sDa9FZsAdqM2Xn9H9HcCV8yRCwaA8pvSO1qr22utcA/kxslO
GOkcsLfNvGW9Hfki2YXujJHOg3xfWubMpor+rtkFiR+7VpmPkRB1RFjbHiRDLJ8k
IVhp/kMUeftFKkndlGLLz1fWGlycOlueN0vrKhheSj/B/ZbajkeDr3eSJSzVOQZd
YT/awrrd+iem9xvm4lJSCRLwSwUErUNXJIuwyvIGPDBOS9LU8IXgLXT/0FKYLPqd
qFBAA5QXeL52VC9v3VQBMgjAR/jQ2q7Qf0JoG6au+pXXx0fmjK8QSnXbOcxeejkT
nHQdR5yBIy18EY8FX3ntQQ5kUzpNJ8n2sUVllt2azCWcdDsY2XuXcpKxp5UTEOmO
wXmXi5CX6jGsToiis5uHnkVdvlScOaviesoexfgXy9L/4YEkR0HaNcfCqHVi04Em
tq8ksIDDlx/QiTRQ8WX1NazuCPaO/FoMqzCamOwsY4xF6S/hWeS5GzXarjpK41st
BqPsidWkWP2o907gwQqli9TcARR3A0AwZhamtUPb1fGp+LjqEF2m7D5iEoYxZYf8
gLQt4e9ZoRfaRvqZ7/G3IEYWVRCL00um7/avR/+lg2CYf94oHErB8aov+B30Kbye
u3OAOWve38UwyESCMeH5gIiIvdrJ9TRusAtXgRO2k4A5iyOAciz/LRUOUJPTyFoi
6cNf++C54pxO/5ZeTju1S5dG4YMjfgjGf/fLJyi96Z4DeBzlW9V1PtDJ2pKmWNPO
qE+xgWW7ZijsQz0ZzYAGL0BI1ZmFKHsRQPXZ6XuVjq1/DiHK69YcDhhcI4G73BA7
SnynLlF3b7LURM0zzwx01wxSP2qekOo9z5fJOyexr9ezJAlshNTq7VDKaPk1bCWk
U9zBPvRx3NUInJPnrWL7cx6LavAqyh7dddlZsTtcpfUs4hh5yOtm8eVpUnMr5sbJ
RuEnOxi5gCvh8svamHwaTxw4OJvQ4sa8FEoIBj+EqXvAObks8QwE8GvqjSp7OeCJ
Zz5K56mv0M6g4LNLo0TGLPlGQXJy24sqfMqO8hZkI7F0vzmLnLDsO02Ioy1ICITK
gtCGVnvs+MCYcjTDQ4YUdYeW9Funh/G6cAP5N9BpkiIA/PPN5rXA45uyQoWm4okX
BKs+B7DidoxP6LoWWYnXRC0jzv5KeifjxCfwk34ZSk5laHdIp6tjYmRtRhKuemC9
BCy5xIu5qJ2RatFu4DsJMOawE9AYluBA7m6u7+mrgYY/M/onPSEpKZv6ZvdfY8/m
i5gCe36Vrbpqa0LV8vcHJX95Q8zUSGBnNaUe1qSpM87VPy3SqfcXXYvjS3DdZBof
uSAZ8q8kfseishFi3JgTQIBGACRUmfUeoxH9rTFL1i898e+EKF2ARQ3txoHY/Ufp
QekR6VlXwPxAkkYeTer+W3b54kW3bz63gdg1EPVJDe01ip2oMC5sqbNQlnRxFyzf
VFM/8QjP+7C9LCd4MqLXjdljx634FZJhbbFB9iftN2mrWBkgCMH2CJfEg5k6VBoD
aV+9Qad42g4HuyBDhLOw4iu286IUiwbscPqQC4ziSDptDcrCddy88yeBE+1FU1gS
wNbfA4HobHV9FTmrw/1H3z32Dmo7RQlpttOluaHrhtfAcEiMuMu3OLyph0D810rz
5NQ7mqHX2LmQ5bF1CXdZYT3Vo2sY4Lxrqi7tosGxBfkOrKol744d6GTOdeTSu2Zx
q927Yx91w8k14Wvt3MSPZYF3VTDHMzTyc5DiDbWnAvd2ITxQNbc+PS5Ri0QJfYVH
lDX1Yv8EUmLcrxKnDnMPLS6TT9CAKnghvE2wIFAOSYiAqCh6W1zQr5wMSpJ2VDTy
QDwT3KsdJiv5pHRSuTPlHcOHaGl3yubOQHVdTn40c5PqY40dwYTOkIRGjhv+FOex
ovqxsZFkQaK/AS9LB/0uFZe8EFvT+fYldbgXppwirMjpct5JzcQtW00KzrkRdhyR
/LwzZq/UBZQS1jCwzGYWDH75rYAqBqWWAZRemObMEsqdq6e1rMuUJy5cp0J7b/mF
isSSb0dlO4GmdFlsnrGgRzLZK3c5NxsqaqLcPTF8AjxQ+8bpi04VzXQ6DLqLFxyU
jjnDtY2V5sjt7i3HHOpcbZiot6OvwB1Se8XGo5h5xr7e99uBvMqzI5f6F1ICD+II
k5lzdGXx0cZ21sSoZzVS1pmi6MxniFMbTqdzHMaRunraUmz2gAdiOlMtJun4fgWW
4DHINq7moWFMUQvCxVLgBy6GAguWh6ahJpVTPBh/Ou2kBse2xmIj9M6cZfZrA8Sn
L1pqfInkeTieeBAknDj2QBcHP06DgTkWtsC8od13SjG8yUt6yPdiXdj/d1heTG9V
1tnoQ4/Z83zviIXdY+BnxsPc7Ht4qUe/F+WV+MVHbg0uE7vbOsy/gqTWgbTC1/wc
yWSyRTBE8NGEMo3OGAGyuetWflJxDanlLdXNWrmjISlpjGoB90qHgkaxIaQxXJWR
NJe0rXkg1y2lVcp4fbpjD4lCL6zzsd1glWZUbfTzr0ehgUNzM9rjEQyoNvXsTx48
hNwQ9mRfr9lDkOH/+eOaJoO/iPKayJ8s7J9Ed4RvURyGmA5iBMsbNVJYy+NBCw4U
p3u16JLKQASW9mTY/lmy4LiaHcRyGomCuA7ohtGseIXoS+VG+R6i1GA11CnH7h/N
Bp5M+K7f/ubEjqhiPC8uX9eOA8XK5RQVSuF+LVUdZX9X6lbZBR3fuTWuKx63fShc
x6bvgIcPwbtFPJxrqDYl0jhAyrefzk9vSKjz4nO3Fp2xWIM+RBPJWEVWD4a0rS5E
CMPoxHDePUDwcqVQvjFGNPvjcNn6t9WilQWD3UvaB5htB8NiGFuPsmTRGFWUEine
0Dy7HaDRzx3A+3ReUcJtMRBUsGWemt23dgH8fzqNQSKCjrYdTeK8YR0r5gFyVFkE
7+GOIQ4ursduaHlB6MfbuK2OpdEwa+jJzge883x9qnsOqC5ZK9diwGFaKVCRMU0I
qNN4J+S1sTruhaOABy7wyBLYPmwdBhmT/4MEtTc2F/zjCfuhUkFxIQ423YStVom+
a054emxSUs80/Qhv3oGCVpZBJ248a2iPTcgBzRfg9ioDBcCb/jrg7oduQV4ZhqCi
80rKZYwqcoj4nqdgqc4XqkYD5j5MRBd3y2GImNGpJXBBMRy3Ip8IeykWnre+Lkx/
DkMFL+ZOi5kd3K4SXZLjZRg1obUu0JnWAbjSzIfYh1M66SXClK8UNn5EgBtStzC4
cBrZw5fXf/XGtrUjAwvD/DX5sZYbWe/e4J2NHQ3pzyVmixz16kLvB0okTmwHX3yM
dRuSzhTcWjDgYoBaSxvrNhtIruLqUPaNjNeiaoXSrcEhz73b4CDvK27quIKlLpjb
AIQaG/oGSaC7KRGulXQ1A3KAJwyzwnK+PFnEZo9qycCI2EYFDh+1fxyIOtfejtHR
g8AP5DkIVSZhts4Aix6FksKyw9L9De1M0WrFSnCIOEsuxiY0+jzs49VbbaTSlfw7
AbkjfNfEPYSiAafkBJtoBnbVouL6S2j/6hqpNDVc7qbZemmMV4amsMW9v2rrK/ho
MxzdAGSVfCz89V4NQE7uBVYKoeSPtsj1iiFgOoZdg2jbt5RK0SWOacT2Wlfh4wol
KLYWuejdNkIULeyGvd73uPO5tlZjU1tuSmjcB5STFeXbe5IXr6RQi3+nLvIuSWMr
CjEa26IBhFKRmwsDENY6MtyXA/G7gZaqQKF4pRHxV/MqHR76bS77BwWiOkFnhsfR
M36a1gGcmu6RmLaMDPAxb97LrLxCNef0qp15pzsee3MpoHzWK9Sq44YjzX13tsTh
mzmRYZX/9P+ruavwwxume63CDCD6H9WFcE53ssd47CkUHhcI+bT8s8kmkW0Slb8s
CEsWqUPxOEp/+jMt7XQqeQRHhbn/RbV7VVSZi34oM2nR5nrS0xqATpzlqQ1k50L4
o9yvWLAG+KKk05/E0xoY+dAncv1d5iuoJbq8X3oc/y1IzPANsfRjFq+4/t/F7QSK
eWXQP3btGAN+TX52k/6lBRGyYXlBKDHVzqjBpBy04neFY+Wl/R4lOjw8vcwx6tgh
OaapAgIyUlKiHydZj3+g3HG9RO0ONvjSXqH5MrU5KkF0H/Gziq0PJIKvRg4LORmH
dtHNWXI17vWpRIbxTuFHaG3205PX1v9f2TH/6rRRzg45hSYaFGUtRU9sxg3UtALH
vlslLWp5eLN60i2lpoFJ8tt7HOGfI0xHknTdgZDNZvSUAYiPzHv9GSpdZHbEXX+q
hlDTPnKqzgmBUMpA4AMnUEhH7c3C8ltSER+Vfz/4jHBHTY3JaEHbiBN8XyfExtNm
hXO3jCqLyg8/iFyS4Tp7IEM+wN6jNx26sAPshkiiHcFdPzCViGtutNDFV+HF72AN
R6zokioM8B4JHLpQIzuYXshsrOUepWkPtsrrbubf5S/OXXLMO3j46AU/5VUI4l6D
17j3O8JnY1vut9u1RRMRfvttHQ4sy39mu77FQo//hjcLTjSyGdq6hDyzR/cQgnxh
p16DWCwk2l203scW91k7aSiZs4HkXgr4JzXKb4+gzO9Y8E2V25ZkCsnHkX6lPIIx
H+vuLvAaEwPxD0RnkBCEL/2jFYchmfBqeqKH3cwDqDz86naZwJn66JUwD+F9mLJX
kfSR9uVgoC4IBSPb177eHCN6CsMzGSg0W1xr1/Q1H04A8OFZnm8HrTIwTTxAFX1i
5qudF1liMHez6/I0Km4bQsf7/cOPBEcWmamoKP+6HpojEGywgRLM8mpQQPVmPi/U
S8zAa+On6+Si30kyMJPHeC5GqboUx+BPc7UGKbdvzNVOxbeFbkuTNU4UGNkV3eyE
LRc/BSzB0Hzlt4e1BFPdl47nhc/mPtLSke2Qx8gb2Crp0V1Y7dYmcxLZxdia9dgd
jGJNDGiKrOlGR6YQgOsnaR8uaYNAqR913LtLtiRYhckmWca6aj++ZcviE21Ddx5y
9brshBPFIH4P6c5kP2OlzzG7n9YIf9VPP5GfIzuCvB06zuD9kcH77oPJlTGaGENM
LHG6ZqbVZJdINMXJ4Kp50v3c4j91UHhkNuxWOQ1Tgy0un65QtI9EY3L2NXk24ynk
iVdRSsSJgFIEsY7Q1zmG1gaeFU431RQn3BskEYHGxk2Dz1Uy/k/FjDoVl7X6G22h
T+KpuBZGvlqHGddi8U82zlszT7pDgPqQU98JLwYu1AeDFrPXWlocNDAJh0SRFmhT
98zHUYGeRmLWXO1W+RA22VoJI7mz97B0/5UtCzkrOpCLe+dgnP6ElrazQN5N4olP
CvYzv5F2TfE2FmN4rgTH2ayDUozLgzsP30IojxeVGoq3ApTWa+QfGYkkdd81Bvf/
i4i0DVYvERV6nYYPy9Gv/alaILKgcSTA/YCFM67U11RnG3rQv5P3zrUGZym0QJQs
cSrwGdJlKHnrRYU/Ao4esdH43EcCNujem4d19ld+ntnw011vP1hPSUG5aA4EvS8G
ZW2kaKKwD9S5bzoVc9Blorg7RHoCzO0i/5LE7/2i/a1nfvy17dELiFxoXXYca7Nv
nvnTk3ncmmZd+TYNMwXqM93pATC2IO5BmZ32CLEPo+ezruACRnkg335qxSqhYy16
/xSzbI6lhd8eVywxLv7/uvBMe5h9wBWLfgjktURvVpYq2jWuhZq5bzZOOHYbDDAU
MseYL8RWk58AaqpsAf+D0lD56iBI1Evh9rBApOAME6eL4D/aB9WGwGJdZsr/Y4zA
BMw0PPcH2G4JFPmlS5FqN5ULjdjyFFD31yBVghisum2DZMHcw2yR+wr4EF0NMYgi
WGx7bNyptw4WMyZE+a1Q2EzDIfBhbUxWWjWRad9r6ot8cQdrozCAG9hD42iKwTV9
QMk585ou1fsPekWPC8C/XZd+njLWQzIKMKUgFD4p9fAcJd9f/x/IFUMrtxtkvivU
MRzE/Ih5M00h878G3tT1Q/6/YUvpyj4NcUMLtzOIBMv3kadOhdyABNf5u/y+QsTX
TzvA2x1ztdwDI9z7SPuGlXz89IO2ujzF09lTu2D3gcZfNGkRrQ6wYx2CLFBXYo/H
dUgC8mX706Rc4aZe8SX9V4GYfo0HCQxdiJ6epMV3JkQ9p+Z4etmK2xQnczx64Fgc
xfszComgkjDRprg7xpMnN5Hz7oLUFf5uREq7x/kfrn64z63ouP1k6blTHvfqcutJ
05Qw5J5mKURNhmnah3upVvVqUQEPJrT9WuKpEifJWvmuCFVfnyu/QOZiD5mfSiJC
aoiC8klfOrFiboE7aUtXoxJGA2Ap4on5FM49N2aw3Fp8G3kR1TgNnbizOK5/4jtK
8TzzLwGP6es7ywOHwTL4xMmjs4UHxWINCMRL37oWaoMVGbBa43KHcBiP8B0Kw5yn
DwEkuWeAest/mI39MSho2N8F08oNL6my9yhxhgQTolsDCOW/UDbn7IcJAKupIL50
b4Pd8a6cQ8Fi8MrIDFUv8bBuQb3WotnCaz4gH4xVnkHzoHZt0VsoEKEytHspcU+z
PEAv60eD2pFlZqWvHFCRge2S4MxHkwS3kxPc+D7h71jSrLq6RBWts6IUD04VFxZa
oWLJ23Ixo6rpTa0kfQ9tuTLS3FnTGor/Fn881Y0PdOt5syiGTFc+jCoEtsjonoX2
xUlt9lSUhYhG4N3IcX9fCJBJm8LfvzetHyx/js+i34ejV9ed4VqhCg/+94SzLn5T
5qqWd8tEDop5fFspcQF0e4pjvQP/nRCjf/LPz/5dfBgBmjNTnGT5D8aNgX/ZbkOg
TYwJYeP2Q9Lxa9L1ABm0fEJkiH8PyoyzzustSMZ28VKnYl7caY4GMy83IdSjtZAo
cvusR1zn/mz7mYnGYE8BNxHtquxRqH1SBEAlyWXkrcSHqAE5RxGJhs6UVXSbkmfR
tDGdOkjHbaZCcuQYqsjj5Vct7tobPRv+hIgf8JPvEiVRwCJbpztNrVdIvrNZHhVs
4TYVGhpQF9t3JAR/KYJczSdyc4ifT1Rg420NpxLLSE2v5ju86wO7dKDm2xt73UDF
HTm8AewVGd+QUbnyV7XIGeSGXkag3SyxoPs4RLj73wiKlGld+RQYmg6jgRknLop/
nkHWlG65vpkodmmBO9A5YvOuQDm2jrW8qEsrFLnodeNtuSJyvq72ZIKHOpCdaVIy
G97WzBG+4ck3ajSq25+nAA+uFPCic/dihR/7XxkTVIaJHUakQBYYJys/x8hpnmmO
JdHDEnQdSV0A/E8aK+Y3tI95pdTIUka/heilaDGQGQLptezkY/vC/ZoGaunoKtyh
y+6AeZEAHhTT1yKVqoQTs0a/k98K1cs/YqzF6QT1tqNSag1aOuhO6p0RiL3jacSg
l6BgtTpJ+4BLLdN+dBBj0y8rYtCEpxqGam61LAh5BOJEE9iG5QW9MC4IwSODI2h1
30k5cy8urI/07RGy7X7q+4xT3gBnr9r3KqxVB3mgwHGBKU0sk6q47g+8jDkEutvw
LAM+dsYlKA0OfgfJTgvuCf7a8LkwD7U1Jm/X/zPU/0bhHThxPACb0WD4cHyxWH/r
VZTlXrTj2BdoYcLVmEwBDL09mZin1tFKqJ8pYSQyTNN64L33pP3a1V8SJ53Mjv4n
scfKmPAtSgELeDLaLJT7PxvIPnMQBRZoC8VCgxpfgsjnAWLNSTV02kDeY/WnAcng
VBBtPrz7DAI1hlsUXqKLzzx07wP4zL2wMpLSjTMwR1jYZhDZqQwGGWMo85dvgFE2
4QVKV8IEXjsQF7hJw6+ZLU7/sNGeMl+ir+aC/ISVDhi/AN6/rZqs3U+oa/R7pcoW
gRPjtzsKSUiqLeezHwIDhzvu0wThIULCpqb1jQbFuQbkkywqJCAkJ3N6DQavyxoH
SF91xYPccYFxuWbcWGgPZca0Me4cBpstzNk+OwoCmC4kijruc5W5UcO6qB7CQnP4
1LK3UMfcTjxqWfVo5rwesFnDxxnMEU457cGrjMl6XzeSMSplGtLer+8kT6K5U48e
JB7s6VQVaDcqoNj3vpfoB8WpBvkUI8kdQMMNQFpTlTAI/qZKrgQmgbvHhCbhuCBq
HU3xKD7Jq90mb7Ry/32xfDu7g1DqHq4NBjPbiToVHdU3ue8fx0jIS7AihPXjwgqf
lQcUxHS8jufy/uIYpDnizxM8z91QA5KNKzYucN3RptmLL0Ye3TkDyUxAJk0JGmJu
9K2V7UafFKnxhynaQqgm+6l1V8PKNj3NoFMJsuHLfX3rmj2hJd55qMEyGY+c5/dN
jTXTVjYwJ0Cr5CjKwNSX2DJ/g9xcjsa5IPyb8Fy4ugExGpID6cO6Q4SmccwQhP6M
scjOMQeo9jhLKa9zaBi/GoRTqOmZ7yOZXtULYKYZDrPczGLQCOygDlvGeYk87fE4
8lSWJNlXjHnHmRXiU4ylm68eu2/sOi1pv+I2KShh1Yek7xlZ+I+bD7Y6Ci78C19I
5DKxB8pVK4rZ/Wl3b0F+NBllcPdJEPoBe0IBKR3sixbtWiJNJZ12Wm5/XnzC4nEm
/Sa6dpCDsi1ran/vG5aA5E/mv9KjG8PRKTNjnQJofI2IGMutqX20pnGsUVMSHD0l
ul0G/wZwdxKwbYAJCiv6OujLRrBjr+QIr5AbZubd3IU5qY2ozJdjKYoBFMJwSpOJ
urlxyDn4V6dhpq7ipY/szCqNycQ6dgts85wi/UkFrN8STuhcRx+OvyUoHDqunDi3
WpoaQp/eDEb1+UyXNdm/Wp/V6APphMgp7jEhPLu9KQRiYrI3ZlH1NjSM+JeTwu7u
aivK6Vv1DX3zN5uVEiF1X/4Z41x6RCy+ildNrs1Us+Zdd0J68s+5L4r7qS+tv8+u
Mym4yKC5NMKAtlVoZvYkp5YgzQpdVVXLKuCc4KQLJqtlwMf3PsI8KcVHpcZigBe5
ClKv3NVpYWnaJI7bAbacLxDfOkN8RcwXRqXy0puVmPFekbaAeOM1URCc/SDOCIAb
Z1dH0ST4fJaZYm0dmTlsZsCKlykOM3Qx6Lx7/HnVutqR9DRSzgYp24UvlGA9is6H
LDdPtp7EmlctcOtnaiAMjdxRvYy8XF4qOFdi4m4EjNTHH6EJsgWdHaGloNc5XPD0
guLuZ0btHEoEdL6rmfcZ5h4Ky28F8J6elSq9Fwlq9RjSKgOoc/xHqvTOzWjuBjNW
WNpT8T0wn63foYB2XXN4/RVcVQAWWoiX4eByQrDCWezGA/1leaT60N2nTooOBgdC
BpZQq2QBfapniQc/g1FBJspsJDqr1EwacGKjTEEkrBqiP3g1pJ2BudDN1VP8AQ1B
ioilV2nx2q1JtI/OLgT8ck4uWBqBEk4SNt7lcpKFufxj+W8pv5odJTnTEFI9Zx6a
P72SwwRLKILdYX8CmcDa2De0blCPyfLeQye09xmkF94gDGqWwgsxGl++5JFnvTAr
P3C0J0PDjSvE0RiMgV1gGcznuExZpx7Sa7dcmOAu0AZLpmDj6sue0EfT2pv0kPB0
1EgM8TcPfUogynRTQsNMAONT6iBcLcqIUdLpJShngD4NJ8nwN7C/eyXnKPzFr80N
uCif3rswXhbnevQSgwqNRFc4FmhxoGKBWbY6x80O55BiQu6NEfDNEDvQMZ1nXMNu
PKmWMl3r704IdY1+wRHTFue0WiZD3Vl8DgkEBgMq1+Zq5g8vX2q1YFQeoSpabLcg
CCTBR1S65u3Ogjy2b+xbDPPFYL/fb/V4yIi7Pp4Jl1V2UWIPMXJEqJVTcpz0UyCC
yvltYFK8PfDVMFPC1q9uFeRy+ZWT5iRSpsPGQCav+hUKRh+oBoO6Dbq/l5zSeIAq
nm5sZ6zZFoRislPWa4Bc9qdLVZlf8Jt1iLafZz9HaHGqMmF+o2ODuxn/hPXy8yb6
fNNKM9WJG0m5DyRH5ywVgqxhPy/WRB5jcX4WVMaPaKv45Stju+yvZE2ariWfJjqc
kt8Vqogcm5s1CdRZ+y/y89M+efbIsI6NyjnqkqqVcyGSE7HwibmrYFjwceZ2J9kF
XbXLDIExqkuFmmTzhnqETnepR/BriHdnjbGx5EMWF5pbcfrGNseFKcwfqjikUMM9
4kCnmYbSVEAT8LLdBGKJlvvR0+5nfctPTQo6F3+dOYm0RsTH2YMte85BJcX+/LR6
PYFR7IJtz00PeN3YD4cGQYAiRz7cktQHlOv63898Gviqhehu+9r9SJyDC3DTD68G
EXRFkwqiBMOHEvWUJqLzf/FLm3FPywXF6Nf1A2kMYGu9fRQ+JiX/x70C30Ip5ngZ
kcgIOpE6L/hUlK62JjFHm+Ksq7IE/6CSV5ZRTpU+5DNJkTJM6jyfYK/zsST+3mwJ
3LU56ty5a/RPT7tXhtde7QDwjmj62oXMCck7QcGgdVWMwHP4KhphM2W7TqFHB3Tx
LOwrUnRHtbjCyFIHl1TwdySX98U7sjTnWKUmA9iwtRf9Jx3X/Kw5NdCQnU+zeYul
CS1GH9BQ8zHxYQcHgFLLJe4O/4p+a6YKmLV/xyF4nsZOAMnadwGt55Av/3+ru0Wg
c/Xoue+nSh+EPwWYrlGjxG7N/PoMPDfG5Rbl/igTZg5mnNk5dEcWK8tmZcybsZ9B
ILrsp/ugjF5dx2izbffPFsoXTw6fqzcPD5DA6TdBRkRUwezFeUCPdXniASboocs8
IKHj6nBzKCvxQUQ0ISR4+a5JOioUQeAYRl0cvf1Cp8tcS5j2Sgg2uqrxFF7p2sSs
hUiuetpD2s37u0c9Qr554fQahrAnIRLSBksZvGfEARLbztb/5rOmgXf5n1OH+2zG
5Eu9tFoEM7RWokCxIDkPUxoeWYoKKQwyK+dOPTB/9NC+FJ8cbnc+v53TKPh9kxMV
KZ2mRkq0Df0E8zb5q0ZSivY98Km4d9+GOShy3ARjxEH5TKnGHUTbiU/sVhCtZVXD
5PgmKwK/7T7K9G+4YoR+pUN2EkNIvw5VfGDBMjbJKMwx/J1o9aFSv5VQG2yNUpIo
VUbW6nOzz7zI18d721wefZX6PDAilKoM78EqRqOtv6pNLR182RoCJ1axjyzgSl8f
2q/cG+hL6MotBgzPKRImSmG77y1Nx6s4TbnwvEW8YafETGqQVbU/BhbEXfwwOJz0
/tsmNXgJfyEN9KHZYMW+wtekujKs4kvvACTEy5+SaJ0q9IYovaQELbgvavZbHlPE
A+lPNmBYWe/4Cgws3l6KIHs479vxd1Zf5SdWt51Q5XRQ59uKgrfrObiWqnbrKFgV
yfj4XZ0KfRVS2GK1GAeBxZCt8rm0S29Arng9U3Eivabi0FKQL4e760qU7lfv8f8w
Eo1yHGzN5ScFpmV2q+2VWXR7xtl2+ucHHPAzSsvI3VkSdh8zrMLXsB+X1DrDTLgj
uOLmg8cO7pbzMNQkidLQWoTll6yYLOYyHpn0l2Nfj2vFD2BsiSZBrIjP52wktSrX
YXhVSHM8Im7uJUYhcJZF67xcECNXrk6W9c63uVrrif6XMmOYv4TS0hDC63I6ygIr
5DHYA1rlFfgucIFOVbq0VTqQC/FuwZDY7OSXLdVX4a9uuGOm+6+Rjgna6nXLkhdt
eFqvqYcGlN8c4knQEqiY0+FKDkwuqSnhDjXpSEReNR8DgDI3eD1hIzMiVmRvG3my
s6SPYk/Xu/B7tswhG4k0sbLDAAqa/65Pk1ppESp/OnyYMXrjgxlVabv4ikRy40K7
w2qCZqyNQSssBceeX9wBrhrvLGwKAyb8TwfKX52QZ5ezS4ItRMWbThoehVytetzx
5AyLTZVJVFousXLhX1u49v8RjQqOCymcmViItkAm919X2uMl2yj4yOGycKZQMmWC
ExOvjdyVFOaV1IDUg6yQtv8V6gvxEqMt+gdQR6BEW5ENOXQ49pvPHiKthgEVTChG
eusakJV4VXxK68724+vo8jXzjIlVGrmBxvp7G1Hs1QCob1Qr52gi+uv7ybVK5Gy3
WD8CJBag1Kq0E2+okEY4DGpdh7Fg19NXuGuHi9BKdchMI9dBuq/m6dVXmw6pNdH4
d6lkdwZV0Tq7/FABrb+wHTbH4SEByEI0xmxhwc9c2LmBMNEVcQkd+wlmO8Kp6gkx
cfVFpGtG6cz8/lMfeBXcpwpIfqHCObs2bN/+4h9bNDcEYMbxtzuo7YVzh6kJhnjG
q93xA3ylgxSrZNApkjb3JF4KIrwM0GtDDtKa6VTC5+r5K0ygQIBkZkhLXb4KusxV
3G23Xbh5fafAA1Ev4ryz1PeFlQcY/CJNv+7qwwCrfVTahA/4wuHrfI4MChjG6jqR
9CwkvpMEB/iSX1P2Je5ZSIye8Dx0OcxHlm67W9OYv6p6KPX70jB4AUwFOu8O6CYR
KbFQeBUHBOQ3k/KvKBdCYdADUtaBaJgHJLrlyZf3pdHbgD4Z/6iP54HJWkeP9xfN
3LY0RORMAwm/d3snR9YeZ+cfhJtGrKL9ZPQoJq9vIKVQBkWXOplIswirA4tXRdFP
NJMQ+hLzmmRnFz9ku9uzdeIRgvu/A6Jt5XobjGJF6lp3yG78NFUbcRyquRC+0QHv
d0XO9R1V5A7e3P66VZrb3s/Soz6mIeDeNbO7wdVpjF4ATyNPdV3m8KoxdUzVj5XF
h3KA87lwDTBuPZAdgcmL2tIFaABgJ/IM/xcDlHq5n2taS0o4Bzno5JCcZ6o94FiN
q5u9AXkRp4JqmhJEhVP0nktiskAt6qjyLe5K1DKrsuhFWkG7YUiylsA37ZHuE3ju
KNll3HfUPXm4C5UJftEBAkQXilLogU+54B70n6BOntLM1ia1/ocM3C4tR4jzGXsS
lKs7UzqP9//Kc6f8H79muRtBqx/pywpfzh+zLUVC5CBqU+S+hQiQFCsgurYjx1w3
dF7eCsyr3FHL5mhgfPZ07T9YJgM+w5D/Bc+FaKJAmTHsLqfCUhRIK1dVEB3t2e09
jlZUIyS57eOLVwMQHqZUKpCrgRHop2MurIck/t9DA1dq6gw3K1VLJJYKja2Rgjsi
HCQwdgFdozfBGbzUR4fc1rIrtDhpnKJh5r8JyAj78CTh3KleGuoi7KwCAEADISPq
E1rYa4Lti/G27sO844+UEBmtKEq7J0mBGdFbDjvEGdo9Pwb2H5aNN4kqh/Z1zyXk
TtPZWVonzeFiQF57ikfCMHC+kq+W4YX4tslibXioayVEPIksWMZv5HW51TVBiVFG
afxnEXc7S4xLyPd4u/2KWrIBwlUghgIr2QRfWRayQ5kGjxQpXdEfhVn29NxbO7bZ
Uo+PLDDOekmQH2l+AiGbYlZ6zHY5W+odthNaRQHHwxc5af/3X58QYg3gDH3ImOAI
sLpiPiG1UGYFBds1x6uXlcQyLa6WI8Aff/O6WjufUr75VQ4Xcn/fhbNsmPkx0BwX
5MWVyUbefdVRCjuCJ5KWE1d4QNSlkKO4DGHaW1iGpXPhCCFdkkapb6ss1cKf5N11
0wyda5JgsT/5wuGxaNrLjin3FGp9SdDTyemtGvuSgR9dnZQOEdMR46h1qHBBoOXn
et282scq5VV/+iUCETKtWlloR6ipQzNbUr2sb+OV/2jL3QKcoBMJ2GuI1PP3YSDg
vMcJwQ1pq+tc9IsnZuuCbOH9TpF7o8euzK95mRN4XP4JyNZcdZavaczmedbF9FoH
QfUY8XWdt/9Z8syy3rRKEFNntuCSzylB5sEEQizpf1j1dTLhEFnaI3Hahpszr4oC
eYfHgBAnQa43DRPZ66qRwwYSQPW/no9Zx4V5IwUPxUvd54OCRPn33rgZXmXORpfg
3a+x4vyfznecWuNzLkrr6Kl+REbgGJEU0YrHm1M3iVgtv2MD1xE+UANGk0pblwyL
5I//b94pplnyxG+hQA5E5KBiIp8sMTUkEvr/JDlv9n6ZyMwEXd+0xYBl0C/cdpax
t1RlQvmAWVhHMO+kXp2EM7FpbkENSZt4FYh/xZsKAZLQKEHezT8SEc11UE8h6Bgp
KflDPlYQ2P3/55ltOl5ydh0C44TFFNLeSOkmTuJGiXF/+fguM27Q7IIP4mihmHZA
cEteZEb6ktj1/NIr2CGammsL0yT8lMM0AOOzHTG4bFSlOl8ozOEyWVZXSq3qZzpP
Sqq8CCk2rrrRcCilOQHx++jGVUpZgy78ojn3wrJftsWzp8D+kLGg6gWRZrKARlor
P6MGACj7e5N3ZRLMF1QIjBgZbDy+du+Em9EhgkKcSvyWir3zLt6ehhbSwLxEFQBf
314JGhY/2T7/8Fn3PL+37GNCa7LgeE8EMvex6j2D+U7C952JtFrMgMbGn0iAD27l
N1zZyWnDFm5CsNrBrWavvCWMkgfalazNfcyd2iK9dwpu7TdKi8Xy0UcRbk3kquQL
DB7llfF0H1u4Fz0OjEBULrlJEcJTxGZN5GcZ3zn/o0aK/6Fxwb1ufTzVrxHldcJJ
JrUagsw4qhco1TAZunYQU2JB8AiaxAMEWlbUbEW7/uAUCbGQG2BnPOVeUrpS3tIZ
eLVBmEWKnt/jL2gYuqOM977miAQh7aPxjCu7BVf5OSYS3+rZ8Sc+RTDu3Np1lNnq
6Y7YtTxJHGDPazraRzLz8xkNjPVT3gec5aBCmWUWH2xcMBimy+bBo3gXumIvicoA
SQVU8mrVRloQ1w0B/USG1zMflZyA/Xxy9hVFX+PZjHrCHpcysPDeo8b8/kaVmgiU
4Lmh+ka3CyJF+KSZ0IBXk5Lf52er+lMC6+Y5Db3UcCZHT5JyIT65MwklU+GT8XOF
M1BjoXQBegBsrDP9hR2FltkbQR3USrH7BZ+u/tWFBppo67cAUL2E+jvLfEhKT1zo
IuJiCrMltz5tYvHLw1eQB/wiN9DgReDdJGTQL05RHsf011jY7sHjb0a1/IzVFEHB
zzysncMsoScp21NuRCoHf8KVl6LssXbyizt9btnNsiRZkh8gW56/9oENIlb3Yj9h
7/dYndmRtqterViMdimOHMzt3/Dtgb8+/9w0z64xw4Gp5gocwkFCV7LHtDRdvmKA
vCOEjsfbkfllZ6BSzBLdTNCe5KYtA6kXixISyqI91Fzr/Mevf+aLz0sdan8Mp/Ln
j8LSdq4YAF8w3yyVMjBrnSlBPr2A/1JHttB/WcXnwoEUaMmi0gNPxwhjkulW5WyE
ja9QRlhOntPYPm13fFbe/IR4DP9NAphK2RWXXe7hrUT3H6xy3NP85k8Jd8sqWgMc
AJi12C9l0NQhdIM1qb9ST5+IU3ljYE/0SsKdciFW9rAy8fhKf9SfpgLKdQ98Ugax
EecqxkZBdNyp2dPkVY/BLD8PUlRi0GEt+gCv9ARMqQkEaAg7TGWOh56LuQ2NMcAa
d4TvzOpVGIqPBTmmiiBhz2PAuROgVkvi377pzWwxwnMwKGMA+/StCMlcVNVKGHg4
RERyZFQI3KMcNw3JeIjMOh9YCwJfEqO2AvjM3xrU1GLEpWVxGk4fNhxo4h35F1R+
PyMiyEjCun33GGQVoP6/Qfpv04/E7G2QHwpsD7DAbFbi2TFYf9HlcH41NxMgS/vo
ABTrS4iL21VOG4WzN6JdEIzrwsB4gOS1tmrUH07STnkdDHHk7um2qaVrJBc1SUyu
jp+zeDQS5yJ9mNXw+9p8EOqUzhCLOOWCVECPL/ardtqhtK7RBMR39IcVUQwv050E
xLlRMiKKcEvmxVIxNACEKEZSQVoZ0XJ79+QJ5OQEAEBGKsE6yWcy4Z/pXXWWRJL/
ZADlQHwQqmWV1dOJXgScSl74PcLvv9DpEEgejAGGjsTjtjEK3353nNjfR6uQtGaT
NdYd9dWyw5fSCUf2CupGGhL9HS+ajs3Nnk1uLDXXE2kR6kgO6fRflaWOG+tlze8Q
q/MsAxTno5BwL2qMLhVJc0yrp5AopoAJ2z6ppWD0wIzzIFJoVOfMTuWwcl6oPhDi
uvpnvbpDdReyD0KjuwLh0rp96RiyTIFOZ+6bqlD1Ia/PaklbVrFc3jWCJ8g27SDo
piaEaT581PtkoBo6rXVjJ7+E4Zvtn0Nix9fvXEvdoKAfHl5sdAl1mYzNAIkdMrPn
qGvK5CmSwFlgj9CyDuv5GfstbOxO6sE/xtGZ4gns0noV6nTwoBkAsXc0185AGPoR
G1VnQo80gRpBgKppSCZZZ6TLgcfGE/byI4xSJbMIKk9oYTIKMXcTUytLqN6yG7NA
1PSoR+kVn5rFp9QiZEegDeIm5REoNnFm0EhBAktgsXpl6m7zH7VdMHiZ5Q1m1pOB
3exAqF/qf4OWcqQTCkNiK0Mij4wZJUif5VPyjBCRhg7Uj5hA+JpgVVzyipsQaW3k
tr0dzjbNJblgC6MuJB5afe7yUHJDzgEbBmwVQwt3h5gYN5lc26BQuWTYpxinEPAn
QVMZYE85OLZ7X1JhMeMwMLfuXFBz4eMfBhneU5L50F+J2wOvg7/CbxFqkls0W9Li
dzvbvsky7E0oHYkXYPhVnbBMLck9+q4FzLZP+7G1CPDdL5zTsQP4oVhHIG990bth
Z932hZl1EklPEXUxl1Vb7gETL7xwKoEn8to9u0BO9h5dDG9t/a/2PZdDO/avO0Wk
5K3LTPVU6YhAsBkS1LUwOx2B7MT0ZHXSUg0TVIgv0M5QqZkNtyLmvwZyPb43GZ4V
cGtwMCIRgxPtB/m7sr9HgyvOdXPl8L6fYhtmZNJm3qXMb9aKZxnZqj1RtuPeeQgO
k7lHkgRLhpiZVAhP8+9gIsk2Ehn5Eq7J2XHJ7NfjDdutmbCFg/qkss+l1hRSjqSP
ewRM3r8HtjBPNMyOnmlBuCeMrVt8YK0gl2ovmcc8j+b//aoxYt8WLAEOsChnD2O9
HGS94F76ESOdlfCtUByII+kbklEX6nxfOg8UEXUDsEPiTr0auIWO4PQLTVNfqF+p
SJPYOV0XU2okmG0iRDqp2+L4J55Dw6AehmFzJtQDFVXbyZGg47K1CmbgWKZsHiUG
Y76qONTMRZijUqwoOnS+zGIZKLXvKf73+9SStQU/KX0lXwcda1WHRq3QtNhRJv5Q
gwPvDIRcHYqhXOkpXQQQC4pYsKCXVSjeDJAuPUz1W3dO0FeNOZH7ZAaSQw4bmXFL
12CDfQSzMkiQonE+kqj5sAqJTY/y05dBanJgjcpbavxieZ7FiWkPghFxspcHOYgg
P3hhA7trZVaseTKdeAg+JwHhXKwHm9dX3qPVn46eCbRMwpE+BK5ARrThvuhdMDUA
Ot37RpmQusQTrcJoEfo0dWMoyTB/lCUVhz6WGXtKQMtocYxWZlf5F5qBXK45tiXY
Anky1MSwZ2E8O/UoKBuwyOMSysG3ZNwObJ5c47r6soU33yNOXe5GTg/VmCVg7qkq
cV0rPejz7jmxoM35OzPN95Wr1yVahg/XzAJj4GF9f9DwPnYnfJbn5nUlsWDrm15M
VJX0Go5SSI2IGPVXUhb1b67+wlavzOSfmf94fel4SL9cvTaMwha2YhEz6ZyUlV4J
7BXVu99Fyxb38z7i9sSZkOt2XL/pgi3q8CBKwzfCxTZyLNZkFOrHVmp+hhvjHd2C
z0hfpGKlZTxUJIFUHme/fTNmARvMox5HNdBz03AgOrunC+izuduPXkEdddPB83mQ
db+ql5blrPJV76Sh6YcAMRZajOFSg//JaXD1FetzlNjJKnrPGMq/PrWvpkYpO+dn
8ouf2WvrE1+zJ4D2qwbSp8/PRrCDML2f8san5iRIctgJpeuEr9W4dZhSGeL6/mxZ
UovJAFEAUVXWNZxZzOCtV41sKLr3qz6zKhrlAiwBlo7eKvqupcJyRfHOVZXn3xHd
SSDKrFbn11NWlS0ihYaoP12+FKT5nXXvnLGR1eaVgGxTNaA+/yqJfEUwL/3SMGPY
y8DorXl5XzqdMS1TGRb2XRcyEdARU3v7gCT+M/2Vl3dE4tjkXv1ZJE/dbwPC+Wrp
EJP6f4ThlDmIKDKksDinsqo3yywPrGresQjEBtkFZzFYAEcHiYIO3TC3Vv66riZq
NvrvFLKAC6kCLAip8PRNUVevY3Oc9Uh+H3qDkcUi5LG78NpgZG8rhBl4SlMU7XGQ
bmZxxZVrZB4dqbI6LhEfJey+ESH6O7SJ1pS79FcP1R80ssTJgsmPgs6Nc56EWcz5
+PLy4INCF1pz4Ys2xfQ7hzevNEWmj6xpKPHA1b/HpBl/RfvZGeLsU+qPD5B8uBm2
BFpdhpu8l1yub8lJH9/xCQk28D6tCOu8ORmQRQBVfm/x2UCD1Tu7VnXoKXBcHIm5
DbsCi+jUO6vO0iMH01ZSZ9t0dgyyU7FnfVeGt+EgpRiw9Bb+/lyf0ADrc3QIOV3i
CmqzXkO6mM56sr7OJerRWZaKU6QhM3pbpy4wDt6Bohq6dJt5jdKMJX4q3MWtOdMm
GzNyOV8XqfdCq3hCp9l7yml7O55zlzHIj3hmKQf4E8SHj3Qks1Mi/1rww2n17yOD
ok6zQrtA2Xqz9Bb0Jrq6talKaKWt6LgjLec+xDlc0cFVuzp72MNHUEnJICvFjtC5
QF3FhXIv18fMahJXEgH+L8PugFTBze1NEbhY+uiqB4yz0DV8z2nWV5qnMhEEVWgn
ooRy165SqGLhyBwa0XdtNjpylkmxTkibW/5UoTcs8VSzT7nP6sJTh2h3cs7HcbdX
62o7OKzjIyh6wSmoC4STUmRc7d+HZoOqYnOYCq73B8uQD/EyhAf2O3wKickRQ+7D
ONlRvUryzTVnLD5mKYgwjNEn8fd1ks7H+LRFH1E3PJ6WJILe01YqxJfX1wK2IJHm
lOAkKY5Kn4DbqRP3Pm7Yb7KddGMra6MG43UC7ILcEbxtwOPkr9GsTGk1gcvNXant
rACs0MKmC0OaD06BBHLR2Ig9mG7hpip8EDayIkalIDhLlXbyTfLWPrXUUYXvdQ+O
GvxFNgDDb0E24AW3Z4NPdV3kI5Bp1KDtK+k7Smznpv9i21GrBKORmO5lJwVCa7De
iTKWzfnVklgxjRoY7HJ1QOloePW3R635nBnvy2jE9ajWRg9RBkuIPUprg6EYB1sb
cUdIA4OYhW0ZV5uwLlmDTmYu1b0oF23fiOFf9iqv0kpeB0DT5GSNizNpQOkxDAve
yifWkGlgGWNslPbOUURyzaIW2sLTvv/jhfSiiADTHYfoGneDC39/doeBOfxNNVlO
6ijelt1s6UcrLe9zfiATHNxVqdaPfVT1y74Od24C89K2l3xNDDwsGgZMOc0L/Egv
kMX40tZNoHZr4LLudzPjUsONWUeKuDcYTWOPmTIlMxQcDj66F/H40UQf/Ti+zmf2
ewbrfsTNw12ZLjR+hgMXeLlahuhRhu7d4OHNIhwivzjoSHOYeif6bulxg0fV7O5X
aObXipKeJx7xNFQWPKBE2hEMy94DQX+7Gizn6lTHAL0zehPqvQayh+eoJiOFS47D
HNlY8j3C3jjeiSMvSkMsrcoXqkFo+NCKDuyncrJpBmXZ757Yd17OUalulLo11Ddn
i/iMW6we5bEPO6NA6vZBqkZc3T9ZCw5MZOsa8dupK87hKPIwCzOPDt8zVWbWs0Xc
Z5IwfJJPYLxNUc+KRM6w1RnUeE5d3S7t6gns04Xo5B8nSi2STmTLyk/0xlMHtbx9
Ia7A48cC/5+45P2Em56WBST+i0jLC4e3sRDyR8RuahP5ZJ1VxSxOpmCdAb08+/JJ
wGieyOmhkeHcsbmvyfGpkNOFgaPuBDVZpjLKCr2oQ9u51i/BthZlopp+JpJhscGa
R6pC0XaIY5BQLkRoqBb/TOJE541V2bZrMhSw6jD3KIIz4vwBBK10XywwQAo+Apt1
40GbFXnGy98AiJc4iCgxNXqUCoM8SFi5KKTk7K0q90cgYtu8ZuqmIj9x4fZRI21d
aq+/dScguP+b9wPzlfOOuSQQsO6YjAyinhr8aMLhmxm/la9FH+kYQ1tm8uqTCsSm
/H6jU5BR58xwQKyqwJW9R+W22atrwY5gkkD4kZSbZNwi9I03fqta2pDQpBuYtp7s
0RaJ9a4IMOSwqu4zv+KB6Y8OEM8ntrz4eVpE09jTCnRY3v37itZQi43e2VYJfRUs
Y8SqQfxN8bOfEG3bt35Ffq5SScIf4yTnaB5gPRSjD5VjaPv7cB+jikFMffPLOwpF
IqJkdg7kRNg8mEqJ4/qdOjQnqjViM7veSebyUegQTAGuqATplpw2yP0A+WWEUt/D
l6Vq7eJiQjHNm9S2V+eiXW94Einq5ynBS0J36uhK+/FZzUQLjO1QBTkJE20cIEnx
1+6QyzagYle/ANhB+vr/QvCT/fnnuXDDWwbYyBizNxjaJwvap0PNfXzl/I/GhkZW
Oh6HbbuBgX2PG+OeBSkW3XqEccfWNceYxH5C1V/FrnRqTP1l1rPmIDFMyYNLvDcL
EPsYx2icQVgw7ArOS8lkT/wiPeBsvYCS2k2NtU73UGJQhktntl6nWKX/lCMpCHCp
iNQnHhHceLGCmrq4Orj+aIAKkOH6ukyriUmtUlBo/tPIz1s6/pJ9ICYEvE2Bi7UO
2NcYNgSfgkr2Lyar1FaEricwtF2tl5rN8DA8X89WeOWcmh2qjnwYW7lz6pLsZWoL
5z3c6GV/AmrGYkv9zJ5X2zzn8JBq6XOqZ4P447JbYlun/cDdWJKvcii/ssPCcktq
t3XGp+e1i8ywJP5icTIhXJxu80q8l8F+wm2NDFguXaGCAqesLz2uoSsHT9B5+JrQ
5qs0c/si2rD9x0vE+5k+j31IHlCcYjuu7S8bMSNCGtFKlldh5aS/20gcoiEPKS2f
S5F/EOwsvsKYGoip6ZeEGuMnSzW+3OMq4aoObZKrQlclkaJWh+q+rTVtnM74Tz+4
qHk02C5LCbBpCVWRHXvmxASlLe1SKrpO5MEIHXDWmTNvXZtNjvRtlQ2zWvsXOIv8
mIdaIWfaO5nanUnb2dE4uRYwOeV0U97FT3DUaNdNabhXZambXmbXPDWL1PEQsUI/
wrei2GDDAnl+4JU1gaFNzcRkyyPSI+KOpo5sTy0gVHn3l6cp7LJPDFbaHi4ngxTJ
8ryxBMwkunIg8UWfPqSq3T5Kek9ywc2IUJIz4HCk70oUZ4QdpvKsmSycvkJZvGuo
dSs+IDMXcyCgtABwxLspGNSpYDszaSjYW+uBvwTrJWC15l/V4j2rKL5u5sKafBVP
4lvwo4waL83Jc/dDipAcgNNmcJb/ZnjFt7+M+e1FEu7Pg0U8Gb7i6wUOF5ZvmeUC
/6pnurhA4E87kXul2VSKhxgVFu8Q9DLsMBD9SwpX6wPblUW9CPJ5eQ1+l32IZic0
LDbtLrSd0i1w2/OwNWFWh8IUyAj0svJWZP7YLTz0EEAg5K56QsbRJot/l7ERTXLT
ex+uAb+Pw2TCGo60HYM9z8Js14JdJr+p80rFv9qmTSisLFmZbuayxiXdFAlJe1pm
16640TNw93NMYmw8vnfafC7ych48KeOGN9tLd7TNwVdAsTs+PM1s8UjUgs4dCUgC
jnwjwOdzOitClfCgyMxcj+bI+nazqqvtC8uqDY6tCN9ohjiz5xtvd7hrWc4rJvpH
rUxzvpq5lNhKPWgpbcwW0bbt0YAvWjsvOYP9xc5STZvl+MAwf0WWK6jnNyrwOyN3
+1vbELeZAeIQFkjGp0wWYL5NG8AWX/8o656vYjNgxqxE7tQhf6M7I5KJAqTxBTPH
ngXIA/HE4trIDCHSwBMSpslDwR3SeHy5cq0GqG3wXaL6dK8QUHpUkIk4d+sgHMk0
ir+otbTmg4e9BuOL4E921ZpQSMi2Tp0sSIBViAtkWD0OW6Sr5rhAmfOAlml8v3fL
SaiM3HFw5J6U/9HuAL84UGabeqWZYZdtBKh12i7bw+Ji9qemhI2tMVfdIucKCfm5
MicyTOx0DqHbRRUUfw+X/rGUnEUY8yo0zZ3BvPJgHlg7kGRH/JFHxbMd7CuibPMM
rL0S7ve7w5OWm76rvG8oXlTc+cwga+nM6DmaVOaFOMq8KPOrnYA3FBliDFzVsVU6
VCqPn+0s97nNM2B8jEg/Lu7DVdDfN8w3AXtjwDwnDHkYhD+QS7x5phjPS3FyXRqU
Zxu0IfcVafL8chVw0bvMZ3j4LKDqTf0uys6pq64dsXLojQTVKV8bYKf+Jzrbz9u5
8RpteWiAtj7+AEFtW9xRObJ0p29675S3O2Saw5BkNBI4L/ikpsdeQP0suZtEpcGZ
r2UeO/GexmZgErRQG55NTB3jVKVxBAG19Ta8qeqdieQ+FMz3z0Sy+EJhsKsjllaL
0QNyMhzncb7uesnDtAInuPO8dGiy3uUA0zxb7YAY5mw+KPyWKMt4Yg7q1seBllPR
wVz2R+9bguoCOzDzd/q4oLJdoEpVpC0qkY1VkZ11jnoTOlzxAVeJqBN54gI4Lohh
wZ5HkN9rNzJU1ZxX9P1miahrrIVXC3Vz4XUF8EGIahwZEcpqFPSg8r0UnAJkcQIa
Jv3UWFW6AVY/q6qJPI3UFZzJRt/+gxowoxPt2EfdVsUFh6/SkvRsTtAUevSRAemp
T9f13RFkXGyCj5HpJOO0QMiQUCxdQT6TfybCm4f18GYdvZR7fODWXRdvrH7m3jWG
4+sYx+aX2q/Wr3suM87neM0QVIs/wOPBsRLsbRzY0CxfvpkVI30XV2qptWPU39+B
NFxsuP6JtkwYSDcbQDUWdG1scsnvZLkT40QwZ+0Y9UFaNUQpemF2iiX+Zz6CG8J+
Ez8kT+JvKYpNzMqGtGXzqnOdYIvOSZwpTqP4XZQAxlveHAMlg5PHB2qmb4aCADM/
Iy8RklRB6udE/zpGTZb418Vf5WVNYnmlqHn82xTGgKP/8GpKTEqpBDB59jTx1KMC
LhdGjRDSiNNQFICBKHSXe+beAK7DZvxlftGYsDwRs4O7wjNlZ6A9DHJ9E6CetmqZ
TeDRapvnfruyFx+MfHMq892OkSBIn2R9bw3JsbskIC6T8vd+44j1oNbL0kKCz8hW
d53dN2PXtxEMdF6sZ43RoDDGCRr+DOo8dwskpnz8+Pfo4tSDg1psu811QmjSJxpL
NOq/bzXeaBgIx01npKfRudU/EUeSUHgn0NK/Q4cQJ7pza0DCoBCFTABeMQ8MdU/l
W8xPBYy/OTusH8EUE9tBv2ngjt3ZjEgRPuN6DkUZIBhZj/4OjK50D32A8F/itwwV
jrSQQtXm6U73Uh2FfZTJLE+1gOYAl48BuBdwm5NPwG2w3J/5hu/JDTUZM3dw9o60
NKtNmeTVhfiPeHIZoqp6SfUFlNOQAs12pT22gkPJowgfLJhSn1EoeB+G/JyH3w+C
VoLpVyZ2JAoVeop4kHljf75N9UdeQc8Q1HQF20yGrRzNxpAM6OEdRxZ3PSDZkh/k
jowZ/xLnjFEV3FZZoSTtgRCN3e1u2VlgOmpr+AzB8tDmQ/8WU9sLnLWjf5WDMzPR
GVKhMsgnG97pzfRMyYvBn1lgCJsZ3cXzKAfHu5ox4/ul9DNrCRv8okIcjyT8eE42
r3ut8qyZi0fg8cyD0AbZy2/fDgebNWVG7D3v+ugkAJgetd/gYBq3b/tS3lgf3EPA
QLBboXay2FcGARbQXm2Fh32j6vCOh7QIOaD3Z+XRr/zmyt9cl+QxvioBuIZrLICg
u0PJJEQSJrWxZhabi+6G5TUdYQ6K6JNq8kUruvmJ3X/W9nN97IlQY2RXxD79J8Yn
7O64B5DBTMNXWBR0DOxx4c6wVhMdWbm2Zoede4dlQ0vLME85DdUi5HMvXHjUUzz1
N/ZjRwvBdCb4VM53HT1mf1uDai/EprcjLeLA0bxd8pBvleG/A/qejmwlf1xg7ZJm
b//DX4OW6YLEUt6VAeYoIBo0JV16zatRGKKfmYEVUdHtsnxFO14e6Z0QlT1WfoO7
bcJEOc+vwc4w95k0gu+llH/r13HTJPNciC3uYS/IZPqqlyVfBy+7hhuUPKTClt0U
9cThH3OiPXgrP9AUtTG+snpMsBF0AyOScS+z+ELW4g4dElwUlh8ykQbOMO4tId6x
8rj8p8sKJcNcBkMXkto1wa6fkOnOeGPtDGr9VYj0bERyzAEeLud7wE1TaF3VyL20
oJnKjWv/kbckFUVLfP4WlnPUTk9qNOjx8cC/kNjQ5lvCyQCBgCxU47bTMH1mdCYL
OfdZnQ5SeP0XrVVIfzYG1KjBfgTZSceKfns+LYTCglSJ5HLP2XB5JsZ2Ax21iaOc
7Y/eAMj+/Zo80TS4f/WPHccx9kMnu0WuoaHAcDuKkEy4gnrlHCwY4uKnlamVgw6S
Rr9mtamfXjQY/PsZHJ1pUoz7ESP3cbdf4vMNiADJXa/40ZyeWY88OQK+4vqPjCU4
T6UoVFhykMqcF/m+kgnLby4yFRkk1e0h/h8MW/zOUVQrm5Vh0+xpSZmBj73zBDC/
bz4lh6qna9YnIKjilpPFyrNPjqKP21UyzrsBjUze+lptvfU9MSN/PXVaWtQfVprm
FyCZUU7S4N4anclpryHEgXDYgKePxxbaGwRdOElJA+cFqBH8qGYuRQ7+831PjfHT
/JviKhCVthCjjhsxvuzAw7BrIINMDqlYwyvrT7MBBrgus/c0tzoIrvNPkndw5tT9
Ud9JVD5H2vqcw+1OVJAf0z1d7H1oINneAxkc9TFct+18JLcuPuWMqCnAz7oiMUku
zcQaHFyMdt+EbU6VuVVhvOpq4yslwbsF65Nruif5HQgJipzUhSaJeVsfHVU7QXrL
qn5O/ZB6XPNRl0+ZIDj1EdTMTNK8GLR5dz0WpZaFIWo9djc4XturBuYYeo7l4LOz
xn6m0OxXTjU7PHBeteIq/ehp8IRLkiMHu5gRAfbT7Q4S08OnJcjFJv+CPmy0egW0
Yx4HHgryyiNgKSy4VUBOr5+WthulRoZeOQQCS333xbgxKJm4JxJ8uOr7drlb36U5
BHrBOS2GumozMAMlZcEH/kye6A8uZvW4CU7E6sXf7tvq4iZGWNTd1elvDwdLf3nc
QnYyvj7hekOCgL09cikNOX0yochopvwITz37FTy91ebJmRkwNoZzXCTNyJw0R8rn
0SQ7uF+9n0hO6eWPYvKdjOOnzjtZU3OZbuu4Yt8fyoBr/R8ZAfh4bihf2F7OWFRZ
znObpcZE0ZgEmD7xehSaJE38sINKa5Xt2pMXUBKqvXG58r8Yf+XKLLGtJaP9H1di
40VKZfWFsjVBNk7TdITIzmawA10+tWZdXKO1hqCS8MnAPlDs4R6Xxu6qKdfMFVmV
FyCuGrN0WvaYtpEYzdUHPnavIAQNQgljHttwGVKZgK4PU5ZfMKdB4Ze3jCgEdKa9
TuLC6eck6MWU9KKdQJw3bOzVv0VWyaSz21SDsA8YoOaX2Cm1n5nsuzjzgYAZwTJ6
jET217yJJH90hXv2F4uB/q7CXJ/KTgabH92R8NfXWod9iqrC6icJWWrVHBLFH489
aI7KuBHJ9P5TD5/1fuY7Mr06zBD860SThN5h73N+0vH4Fw4d7Roa2DCHhowOF6CD
OxQQ9gQFx3Tid7pTVG08D3hEDw0CHd7C3p01w4r98g+XIe+62Qp9UiO8kkjRPfIx
nO2MKueVPq+BlLmpyst+s1x/gV+uCX2m1BYsdxmIjDyZwK5euMWXF3EBXt9ABl87
QYt9rlQYXuLpAH+UhIG1ggfF+NAcyZfuGFPofAlMHW8vlddRRxaQaQ/e6RI6O5um
m4ViLYlsYNHSQ1KwnaGYK7PTD8aERv2Gj0SGZPyUfg1id+xKSXNWkCswLVOz0K06
YWOx5Gw/BITIqSYZPWxfnmDA7nNq7URUZfvrJtmgSm2kpFoxUziKt7MfSHcX+N08
mQaC04+koxz6tgtNDtvP7JARqMAgp+k20joYeYqQc7k4dsiZmTOGDpvHcRh5J8o2
FdxSR+3pXlMPlO8bWteCq1P2KcGEkPCsx8YXw/h2XKrIeCYznbXmlwrOSjrbES+7
bxIQyrBVIjXasrGIYGAC9vSUyUoNVcZ45nnujB3nCi7DBmmfk32BFongUU/T4ugy
2TtsC/R8O4bG9b6HG/X8mlfa8uA5t8VLOhFErO0iroI15SLrW62d9D9ZoFH4dvr2
NuUUZuUgHsNRpOjI0tAr13cRJC4GMpXW4ZacEH8jHuMuvZ6s1qCjYPCNVbYvAoBk
K2uL5/I4804pp1jgRBHPCoxV6aYdm4oul/HPPJnq65LsFNungBzfeLdIPWOteW3Z
AmFtNDuZ8l3rWeYxMjAUnFZ3WZNfmQ7QjjV64JLECdNxQieOD40DhHKG7DuuDAGv
s3m/WzfL74ZdPf1kpBjXNpXeo3vX6Pa6gWfMc+qZ7Ft+ynge36TnCmADhpU9fa53
08KtOE840b81uuRykGD0m2Xj2dJrnmACpxjfN4hvjdFfA6zBFfxT2DvtOcBdcLiX
d47JOyEAlGhPyql7wh+TgGX1D1rKwVM78HagGyljfIy0w6GYajGX6DaYIGLzYdg3
orIw0BfUkbNv3xKGN4jADNuL9WPL1FWpEOzRndhEjkzfK2lBjsO+u/Do8VZsKPop
AM6owt7Lm+P3pc8v+OCtGVXUqEQxowz399Xh6p7JPDMtRuBnS/ByNbBaiWoT94qk
Cn+zJPXAJhGWWDEsW4CQLiubLAaE9gsfkqax2vIe2lfX67oiY6rRhBd4eFxlR4K1
78++W4ybINsHzdtaCiERICOhYPK4V2gSPyfMhG8AUA+ZB+jMllutPHjqLEpcFaEH
ozsjL2a+h1Uf9utrRrg08VXsuwn7L7DYmW8QMJLPqmSH4Cveo8BdgtVasYg3assT
DG+U0vHNMbiOIZByhVSCcJ66VccCX0wF874KGhxY+08YG4xmZStgbG80x7yA58Sg
deZKB2S4TBF06mu3ZF3mAnPZiiI9dhZ8I1+F826WfiypQ3pLkqU7IydSBfvtEjmE
GZHVfTQjDZLBGhd2fObJykNc46B8YLDC7sB1J71b5J/vLZniv6KMToQ0B+7hqRzV
SO3/v1r8fYjKjrwIjybD6bsUZrsy6i/yH6eQHncAcStwunK06C5Y7sngmdKJzRO3
3G+yYaSZLcgNfZSbp6y0TZiDQjarLVdA6nwl7xSuid5NjeIaiuCTefHkD13UvbcJ
Bz6OcuBLCNBS2602/GdYDivMY0SoHyH2IHMgwKYLo86JVPUJGa1aCmba7zROOk9/
XXRYNWU23sAtlhLyEC9yxS76vMoK1CVnxixDFTFYI8J59GGJDJjqHIwU3ahSnjWx
qjOl2WaA6c/eOS3dVEvX218rsrxjQ5Q09GbibNYGxld/7y/otsoFnQOIEnG5G9lM
IU9EbbQojpwFbaWlXpSzVefr8a77XmQuA2nFRTYFZ7fblrw+Y/bkrdIkzGaid4RI
YdTOdk98Wc9rJkekpvsoed6CyBAgMo+JTpy7iJw0YffrK1M2cj+b1Ez/2lYnLGin
AHgRhSxTdJInUtIHxUPfcEsOdW9++ERyb/u2XOXfaAW9k5pbrYKrgn1yiJD8CgxC
GEFNq+06k/u3b5Lui59EoAIt98i3z0U8uGJisth3V2GYatNp8n3A4Ik/Xrndd11z
N3JKuCmm2fjJKYmhVGKbnlf6OL4oXOjJx3vmHVwu1r9MV4pd6yk39DNGxZ3xY2Ql
mnyiX7UovRvoGoabTT7LeOE3whLc5PrcnmW2ZUf3n8EPBMBb6V5+JSwmUHuWapfx
O8bLC3Rf0LQX7lfgD3IGRO3DqwzyqZzhuH3O2aa8jcnZK0bgCJ0KSYCMc0UF6ANU
LXZSMN051gSjw/EtOrokpwr1ZEi83AQPgh4SLylN79bDwZk9NM99JCx1OgkVAmlu
Mv/s7HKjmscLUVUDeJYw399ZEtNXUxHxss9ChF7pCUMMvV4DT2PGyyxbxtZdDi6I
lhMBYU++nv2guDtm3ssBdZ/xo4G4Ls8WY3wmWL2+nGYvU12qLSo27AFEol4p1PzB
gCo9GrJ0V/NRtzzLSzff/KaUkMaHOABVy8V5yxF1lNL7/rMBFeEoexxAbQQfe9IC
9zSuAMp321XiLsa41oXtg0knatHyVmBiqFmWBzFI/G7a8lGY4KiRYuY6rkQ44k72
8vVHdhsXWHBt09a8Vw0WODjYb2Xx38WGJ4+ZYUy2OcRpGiaeCbNmxsNd3yuH457v
3jCUU1CeukNdGlWNuMdRak+FIIm9QtsMHFET230saH5gw/x8HWNVI5Dv8eGVBcRt
u8OqIWxQdoMDFZsfPOyCACaLIYiI2p+f8+mZ34AGQp6dg8JoWH8dhYsdcCmxUYFG
XkhSe744x78PR2FS6qmlkAj06rYbl5BW7YNOvJXEYQrfIX1tO49b+Mh8J4sOeFqt
4cXhLvVTHku8EWR5hSEmHHWRGKUSWDF9BmSIkpvSZjZUuZMM/kBM1gata05LxV1Q
+sKcE6JysytOzWUi8R2/gdH3gJi9TtDWcs0b5QBQHtIQPHfR14mPYWN6UmE6IaC2
nmsp8LOTNqBbjvdHBF9TvyBZTosYMTy8s4qHqh8kFvxaTHMugCU/F1N2fDakIy9C
PAduvjZXYkywzzOaym26VnidhD9483sj5AoQQKYN7TFwHKtkXLhy5ypX6/3oNXak
vttOfJHuYja+iHHrUjKnWgTZ7JRYcNteIhXpmBtemvnqU47/f3EpjtENNgBDAc3L
ISmjPwoz324aa4zizC/3Yqjai2pqHIQBrS1znlT/h2nPlfNQebP0iIHpeokF3Xis
ZK8ZeHvy8gTsxLLXfrQpOPM/Itaovyjd4ZvXxLL++DVlabURRjHvtmMpT+aoc6zk
CWVGoKkgZWNAXP1GHqnUCKXPbXHhlIqbkMO9HDd1/Mq6P3Fxxkg+ae5EqtHzc1ON
vscwA0cikoHfp6fE9yC5dNOrDf8upigM7aNzguk2olZKngvrJhWoHpUTYVDfIpyC
CevffPWllKNyrGvgolUrGgzQvjUF1PnGfgZb03ZoWDQy1uqWpZixARVQflyD3JSK
Oa5itokg0a75lo2nunvroyxEfic/239J+SyAR9E0taCIgv4kCxv2Ia7F/zwytaWu
E79lRCwEWAmoTXiGbIJk4NP+BNBdBNYH3NdsxZiQMNKsLfwn7Q/BaAhHpuD6Y9C6
zK1B/bImNICWmuEHAh9FkgEVK8NvSsAQJfeGvYlS6Qrf5k9R1XX1GtP65apKMBsc
UlR2S0vil3cp1P2gPxc+u09cBCp4dpNrtnV5Licl0aHwFZ0aZCU9ZngnBG7Rs124
dOC514sxSRLEp4qabAwCNDI4ZNm7iG9C0ZtC5eF49wZaLgclSs47GLfxVBtXe92t
vvcG+cLuNldQQijZpcvi9LrsEcentuT2WUFusXEA7UMwgfjXFS50U9JuzDJK2e/d
9kA6VgRq4z/Dnbh0qNH3SMaLf32M+mWHD0E6vqcqEpMvsag2NJoqdxSiPJ8pFqkR
WPcHXXpiGhruxuG6ufTDHdRabss7f3ovl8AF39kQktnzVKsfxgwoLf1fw5mzY2sT
UiUN3ceGEw0ask7XkqBUzG6nScEkgIqRdQ9vGHO3ebFE05qpQnbTifvSn6jzudg1
y6vE8PnVC3Ydm+PaT6bLjXuvO/mw+iIQ01eMZMWNIjPAWxaLN/6fkKfjbx+Ga+N4
q779IFFN/wUqsbY/rchuPUJCSXpDup6cuYQNduQjEoPvryUwhHZqiXPLk2BJNIcA
9SMw/Yz7uNsp1tsNmlp6p7AnFTnRWQDmu4YsJduTBF5mRJ8SSDMshyqCb4u8pEEE
F5xBMPRHdx6mNm/x/ua63PoNF0WY7bOEy5d9mmFdhDgo0PU0pcQTiByLLCgOCgut
SRiU+sQs9+nVmREa5EPzFPGST7MFZaXw8ob023lgv+27A6dwnrf3L/ot91doGkmU
C+nzLgZNkdMiYNGkcRasgswF1fuDINaakY8vN7nJpuL3SQnLij+TdqOh6QLkzUQL
PQ3BacCNQVRhsxJewKDVsujeHS0S8U1OdT7AsGrqvu7LI7BjXBhEO5Ds/cAtsqZ/
/REvc3sbEaB14BnnZSCWGK+T4kgkKZK16ZcN/zAFXWFjcZv/aqmUKatqvAgaJsA4
kFefHnO6EnoiCRt/REv23e0vI5nOij0v8Js7Ulq3ZLKt05WpwS1JkD46KeAx19Tt
JngrKEkcEfAVlQqLSFkqxDBnh0tNXjQJlE4c3Luep5dl1Vbgm8tWgWPDlPE7q1Ko
f7noIVc7j4rQi1XVfD89k6CAJHzemtojJylbfmNHQxAvgkpO1vdSRont4xsCT4Xa
UcLxtQXgh8WgUbqgGSPcZYlIO8xVFata0YCSn4arvdKIMXiaUQuyrNSbDk+btPYV
Cz6y9rWrFItJeQ6yZDOkxABiFSMZvuKg0HyiTQmzpuQriRm/KL47roIxt7wPUNpp
5KBjNtB11rV8U/i3V7/i7rWp/LYNv0i5WFDjt9b4pofTVB3BzAy6sAmjV4oehT7s
InlCfAoNVX5dmDZ/KiuiEbmdudH1qrtm9EoYw+uB251xwND0ZYOPcqMRRhuL9arm
jKftjpYB/piTp1347myKc0aWjgDx3BXGnptbeAznCc0IGbeNqIn9wYSqlOXuG9qG
sGNPWJKiL+vWMxh0jj6gvZi+WbvyImuQ1g9TwWerV4Kv7azxmppuGIOuubLJaA7L
mB5lmfKNrSom79Tv88sDFlkwz9wer8sVa5qWRUl/Sosj39HJB87uVtNjcqk1i0gx
5j4iOLFrp2cjG9Jx802hkhMGGqIcb1D7prGOlp5bGz01pgOBa0+CLY6kTsfcAKjH
bUfd03QRkGNDXaYhDcQ+G/xWyTeqOKW8QhvqNOHS35oT2/ktEcLMMzyhC+vMEsvU
qge/c17D1V5mXu9NamxicUSMymX5xlWV69UXTKI7Lk7c7BwvmHN644x8WFe+EY6E
TdwUD+PjhxujGrO/MV3QmHP2d1OXszKHhAAqEzPQcuWyeP6scjSD8NyuPVPyXlgr
01McULGc4vRmlO+A5VdDTzQBHbcFhBZ1FuK23Gc4nyiR0I1qQHHj3mOvSIO5Ogeg
6iwpXjXOehGq5LEaozaWQFFQVk5hXMFIgBIGzgA3sRR6z/hbFYbkQVn+09ZmP+if
MIClVNfKVluI2ofrSnzxGWQZKCO1jFhtiR/QVh1aisEQKWzsR3A/BXNauCvskLlZ
4ZifviEmdT7XamGOFdu/szcRQIog2Buqp19IILVCBp6AXSAv8kKofSs5E13hQguh
s2ajgRUb21AtBFknZAkaIbiab0JJO8sYVp+UeGNjKW33RytCGTxt1oI2gMlMAlT2
r9Nmo0QHXGDXE2+z/lyj7Plp6eeKGaR8yWIdzVGoYolceXanEhmvPc7wc3W2AD9N
9qgwoZZnNh/fWUJ84kbPl212d6dEgQB2vobV3HFvOiz/xH3YFY7YSIs0Yhps1hi3
O4mulywliDe8mOZ3bQfNXCSW6TdBkEYwigde2k/tyqfVUCbeSxwugxON2bA4iL5A
hHlXkb3jUCwuowhLWi3nqZdm/CIUutQOVAtEIpeQmbqus171XcCjRkFhpg4FXS9k
zrmWA6nApd54Y6lCDUmpU1deKBZJeVNQxfBXAoRCs8bsJ7Sm9xSLXppMTwwY3EQU
pdnewg0SSDm7ttsC24/hgnPADh8ocqmgm9RIZ0Jj80UJ4MmntMVfx5LBKtdpl2++
jL9SRsDQ2rf0Cch9dv5Gsjy75lDy1/uT2rtrKzyHcFPv5hZAc3JOacMWBJMTkOUF
LRW+RcqtlzKgyHabu8qiyzd6z8aGYsrIN8ogaKEZvZvsi3hRNFJej15f2WxzgkoT
NtijAEDA08/KsHe4POQ2G7RmFAydh8pw+ElC7i3PwcfJ9vg1jcM3J4+XdjDjQU9P
gj3mVxR5wvIBjW+Co30+zgP5SUP2/SbGpNSAyjizMK62vHom6k9LWXjiqdzoAFJo
IiegMKjWWiUHbOERysXGqqI1qVz9S4beKcZddUG8gmUMedoXU0yhDR1MslKyXkBc
bERY8bGioUG3un1zN+WAej4Ytfp/PJ8ja/3DkN78HHTyxxJEKai6PUGb8IKssD/A
oHMBgX+of+je/1cwURh9CwCMUXtviDVovUIAqeU4MiYZjlxIx26WMpZTy7Zms4+q
q81B9pw/nw5D5qnvgv11MpvVaYgbsKq20awIsoODryvg6+H45sChAf8OYd32gN03
9XLPQO3pbxdieYl/MdoYqZ+clyHfx45vbLMA0KriYa9jalz29A2XfKbj94I9NQwd
YkDiH8DNlyKtFKUwOOR7RxIHhZgNmLA3ksOGPc2FZA+K2JIWYNzAdXvWWJxvdysY
7uhaoBLUs1FcCC3M7t6LHpJIFWemDmQZ8rFAJ9KFyhr8GArE0kY2S1frm53DGmDv
yMPB1tf+A6qHJOUvMO9kdWOKOnwX6oFwCshM07nGahVB6Kk4vxVrQG/sxtYLL5xh
xmJ4gZRZbZACfbGjIPhKxZaYvprLXzsruuVC0AnUsxtWC4bVIOCQ85J3AncGryq3
vHcsSiUHnb5KpOInls7J/DTiTNCAWGs+LRFrP7KXAq/5RyYN7F80TmBh/FKsBS4Q
v70RuW68RNt2Zo8Le5koIsi12vDDJTHZcpz+W5Op51bWKQ0P4QflmJsfGN7pxYnW
Vi0oXkyVhpPIUBmh1PIT/d3EgYWhQPKH611gMilG5lWfdlCWgiqAA2yaTxG/zMJg
yfKFhdY3d/WoKvC8fGPXM4clWvUJTiw192q/osPLnuP2dUFuO58enuHzcc/cJZVU
ioMPPVmBicSmEkFykrHmlUH0bwaEttpG5dmnp6WwrrzaPFQYRVuORSIV8ockdIzl
RvSxVoiK/6TCqc7/fpPi8V53Jn9NykXEk+gMcUAxJ4nZ7bQK1jlVjUxKqGoUDTnM
JZEIRPsgRGWeIoyReldIHS/SsuTj5Vb4K4CqbTxjjJ0i25kpc7Cl+rkUW8fs0oSR
WxkLQN6uu5wPcD/RkmpqbNOXuaeSkMLSdY5AVlGqn2TvmV0liJ/PosUpaOpfHLpH
tlYH1GJ9aDIdfFy6KUA0GD1lOEHz2+6eY49jtoq2xNI477+RLTZLqM6q3YlJam+e
QoFa4yWqDlH1ABc+cTsyJyAYhwQBt3QUpZ7naW1QzCPIKLYjC57uHtqzkVndWWQD
NFS+Bf3N9FZOY1uzmwFCO8EzGgKWYE3NwvusWBitmHdXLyeDCLutd2HvoGxxYbPL
twSvrdAxyiX5JFniJwNGFUADkH8SwsoO8U59duImxfSsHyWJmmRlIgaiGA+Y3zxW
Fnw64i0lR8OrJd5crYzVoKRrZB7QPw7DJHCO8BsKjWtL4BoPQH6BH2v2bjxL5abS
W87/QSYFyz/oqP8yEcsl4lFz/YzTQTFkul7oC0HqdjH3MQK8nGmrDWnRF2Z95lIF
SSqGVX9aqr6oYzQ7LuT/Z5pDK0/1zsu8rwy4stWDyyRIYik88uC5a5tatm+8LMfo
k6H29dtfV3FXPzNWCC+PC94JhAqIFZCbnYsEvHSasj3wagkxe+A0HbN9eAUivN4P
GhwpomQ/VgFSZMabCsxSHmhomjq89sAY8YrDp13FdbkjUl38BR+jMmTC5P6XgaUE
hMVgN3Rp4I7+ANx0OjWFkM8b5zW8kgrKFtihcQQID1dRK3z5iyB1/aQYL5izPyww
1kBCJHMzDtIzyokcJa4LQWvXDSn00/TOqdrCL/CubgNaPJgpSoN5K6iEQ91Yk4vA
uv6OakWHzoulabKxa+iytTAQHk6ArgaTBEEdV3/HPeHlU//O9GtFFE65BRnxirbD
h4HZx/RMFFti16e1alUuUs/DKtDxAPKUZh+lU8isvVIJqh5sWezaAOj50cbrvE3j
4yqvhYni0akiSigpYwmfstVjKxcUersh2+Jkt5R/GYfFsBlVR6TzglgUoiKV5Dz5
D9YGdP8PQDIPQkv4zwMvP4whceaDztSxml89X7uX97DPhdPwmOLZrOKZK7A73TdH
FF9cnP0TVszwv1u1fBkY8ICu8Q9qKrho7F7sqqTHA3bfV97lH/bDRPxfjaUPq1Xm
RFvAtqj/kBb3GGZtEsJatR94Z5jPVAIUKyge+GkHKKFA6Qn/n496x3fNWWRgNQm4
Ep5WqboI95Sbr2HWlzJb+vb7lfvv6bDUba35h3pv8hLTYFdJoaNauZhlWSFiU5jB
PaVFDIpzdhey92GNul2201ZTg6U3mDbJ+zokRstfeXGKkZkm79yi2iGvjcqUmix6
t8lDm0fRjIH4PEKXcjpfzQYtf8DneGQvevVLuj1VATTGe/DI550FgL0Nn+ERB4YI
sigPiKXocYsnAdH/nrTyq54GjKPh6T0gIG36FTfcZuxreStUzm08QdqslUflCm0H
CCBXw3B1v2eM3EwSySpt0PYVaoLKk87LJwFQAYY6AdFGblMJNH70aMCb78bIcHaW
4uVJ8X3pZpy1jvr9jfOxcr5o445caDKvFvHGZiqfAVhVCrNKlocSG8IttjVV7F2q
IfC5h8IWiNV5vkuhXSvLy+URgolk1WdqBepiK8CsoqU1uWvvkEgt1tNij+6C7uYi
b1RKic3qnJT86gofYcrzUaTiv9F+aI2+3Sigh3Xs7JEmDEWqz4wA0X7dKQoBaXQ8
7LXPpCq/y45Z+mMny6bgxVuSF3g8d++o0gBtgt/pci5HWzMfT2smnM2UA2ojeEGK
lLoLHNT+F8m2H8AxvsscJZckmltuosEwt+IwjzBSLfUZuEjY6Bs7Pss+tpTp9+Qy
sFe6tg/kgdJNiqP2s/oULmAVXj4hB7pY5aTfdoqWaepJ9inYbVSSuKxaMerBu4rq
nGX+968cZcfRdOp9KUJRxkrB/7GLb9g4DQziCCs/4qtW3Ob8HwvHPBTCI6PqX+zA
5dJ2onBfV6nfgCPOw6JN/RPI/E1xHsxidiYqbnqhTdxotBr4Zr16pRASE9gmHjHD
+yFknE2LoZ/aGdBL6mvnTcL3MANjeq47T20Ed49QTlMHcBBjfHnfMzPHePjI2MXB
LydktL2x+hSDUJSj2BIP2q87CmnDLKaqU2SA5Lg3ZiX0DoSEIxqrDnrBRs3KV4zx
u536svKdwmIyKKjpoJ7NF+6v3N0wxCsVtkh65QY1MPut0wHp2GOZGinRpIcI/qbg
5n546z5VNpvc5qZiXiZxaXJy3B5v5t+QmVjV6VVjGJTcYZ148fAVwIVeZCDwMFE3
6/Lc0abPXh8OBtPxCZ5m0d+R5vNlZFijxPrKovc7x1c6umtgfXTW0XTwADwxgjnb
7GDwDJkq/JKY2OfeejS936CYNUv8deguctRur1L/aR5i30sXExztN1xHOChHpmFR
ZKA0lwEK9HmMksKfRDqyTmW7eTkmQlTBiU5MQOClnd/llIYf8EdXh/Ouoxz5EArY
PaV+m2PGMR8BKuRBkxaAxIxcuCD6kuCayh7ZPyi9VC2NiMjENjhM7OJ7ap+D8cu2
CQQYMAUIT5lqzfyTB0ocHfUYLa+D5itT/R2a0B/xGlRg6eQr1x5OMb8+PbaGyZ0N
gANTX308jMS0H9AM8HH18RTVhHThPOtVhXY4v1FnYKRf1Kmy6rPnydkjLrF7iEWl
s/ZRgJLz2yYCj7jj/LJ9X9ErQKqh5608V4HeT+Nvl75l0G/SfKcxrLA26kkeiE0G
09wv89WQF6wLZJIt+fo0pcIbm4J5wwL1G5lIR+bwnjsbqApKTgSShLlBW8iUvWco
QXu+MO4LqV5w8t0NCiK6IJCIB/JrxynIFZ1z2T+jR4wDeF/dJyv33WXt4ePrprKX
VzyoLnrhClNtIwih8xI47HOWvp1u76TPcIrE5AePUoaJuNns+0nYbjWOmhlqqeK5
JQMF4zSP+HPTWvWXtuESlTehC4W1nhiFLBCDqIRjcGqfoUExq7R0xWEhoUQZU2rY
BIkEZZw3X6VTL8NtgFMhHIL1WNYXWXv1TsUtdjj7UvkBKNvhZHuJaROFDXDpXFBd
LXBbgDe+qIxYFMv90GLHpFZOlLR8xrx6x7o178TUCQ/ihqvpYYkTbc2JHqmkV67m
XXIGoFzCnzJgisDmJuxV4SmkJ+aTboHMivnBF1ngNbQiu/JpLMoKxg5xgtFefjN8
wukEKXyjseWg6IiXf4r4ZSrPbHNaNBxMMmF9D0lt1LhuWAZuFPYxw8tebG0lRp/j
Nm33RqLEn/9XBRc9+2s5AiuqBcwBklvGGCbUD0nx9oTTUIGqRgJPFlmP9gOiXiRY
pkgtgbovsHKRlm56vlvqLVeayVwXuSgDMG4inSLHydHmVL+njtGcBdiBRo6mBAzl
tE0Q8ai4Kw8VVwrLHLhQH78P5C2zXkKMrfw0kxWQogkOU8y7tTbcxaWc2+8RShEc
XaPkViHj7jqFCcRT+NpMqj42IY41qoyxfbDkz028o07SbQ1ACJ0Muqj4X3yNb4He
dz/I8+gbKb7b3GgPn1Px55lOOKXzB+caWcNU+IYncJtsZVucUBADmabIEfmKdJ5f
w974bBxn85jgWGr5lPurZFtX3XEPyDjYrvgQv6pYV0carWsI7AbboDbRrXZvWDcl
mqzGZPiKtMZQralVLwJRZiV+J+iAwaSd+CBOY39YXOcd/LMJ6wsvW0cKy+mxNZ5L
Zx6bc9UWUYVPRS7JG24Y+O6+hIvaswUxhs5p+FJ1gzvBE+Q1JQtxX6Djx/E16IIg
kXu1YwpKbk73XhANZMTBgu7amTuozuwT/gip68v4OGrV69+M+quhpBe5OPRaEc8L
OPyix4I9/eGRlRH4+eJ3ptIksZwRyel+/cE+A2oYR0LTUxd3NtwSv7yAf2rnDtYz
j036dvwh55UB4G5gcYecQJn18IlThS8kgpktWmedm8lHbJYw6j5cbSGsEThMK+6C
Nq0T4KByFDqU+JaPTf1Zj/pseEneIaI2N/D0Y3giJCthr/+k+UVA6DG0rtUglyHP
UgoiXqGPEYd9TTpb4iEoDpc16hhTo6A/h5znBcewnAinJs6YoGijIwm7W5E09gCi
qDvaRmPEEWo98koD7T0tNkvF3CgiBZBSAvOtqs8S0bQt6O3imh5EXTJAExTaizVM
GzG2K5jt2xxAHNIoWrkuf7qdhfxnipMbodGf1fUbCBEun8HbTvnQ1olZSjyQfcuS
mrOPu1Ojq0b9usrAFH6k6hKEvngLUD18ESsTBKmzv7LQZRG2gfwTCeckp+xqN6jn
PtWIx8PdFzPq1LyjWV1MOwvPMDx5od7xE52fXTbzzaeTUzIGDbmP7x6BM7lJIu4v
wEkpklg+uY/TboyqRnuciSK2xm1727EnaneCaXdoandlG//9pSeYjRGR/gX2lns5
ORUM6V12e8fXhOUtAWW/JoSjmshlGzAe6rWY6rVxwQhcohQbdZ2fg9Ubf13c+yts
4Jlc4nWhkBt7Wht23LdrZ/MobkDWeRf9/Lo9PqA8wi2VnFlZgpeAqN3w5T3zR0V4
T32G62YyBXkheo12J7LB+R1+QzQ5PdTeaL5oj+MjbGzsEoGA9Cj4gEan9HPwg0U3
Aw5tX36w/yvPQPYtH3BtO2kaqima8f3e2Lxw0t/9cv8V9i7jTtYOWwZJ8gvV7vfz
eFPqTG4m5HecuVLde3FTXN2f1vf9BGC4lhk087ZKTGPs7gaIRz56k1DSLv34Jjwx
E3M9z3ydO4/Pw4xQddjCXHx1pjMFGJVvE6pAJvqMFQkLMxTrHAsHyAkEmZq5O6g9
XqEJ3kiQaXonUCMoG8AobDKF5KTdctCDnaTlfafqJDM3in/WI5z6TPUP0d35pNus
SOVpGAf6j0xjII+PBbkxa0BavrpyK5XGhiOm9OJdWpy5Rll++bh3vaSYjwqTGqDd
YruiRWF7K4gsualHOHAEMmnKt1DJ0bY2Rb5ehiUHX/JHfstyXMZ3OIYspBMyuczM
GQjS1oSHTdSHkSejSaKRg31AddzDQbb1lFetRAwA6Eo+GWrTvKzVZIMpBJ7wMd9T
8TRHfKfdL5WQiCleJMlRDmHhns75K/rhvhh4FSJKy4oLIlblVBDELFbBjyFf9JjV
Dfl3kwmfmf3cgAMICxUJ8qVXOvtt3Qhz8j55TeEjsDxfCjt1PllbsbAUbELTaZ0q
E79MTOjF3zD7AZzRyp6huzUaJJG+2Q76VrC/k0UB55oRTcOgv+i3GUBr5cx1NnEo
maT3bo8pfoKJb0gftuqW/p48hmqTUHl6F/56Zu81Z/M4qd3ccO6silfB7ciU65n+
UxDIXOieAY7AsMHh3AOuxg64501II5Ngt2pi44x6qmCgekFfllhHFLUsEL/jGIiW
XRa0W8TucSDFu1/4w0/70EZAkKXjs6YuOoy76HGgfxpggpnIlWgaWL0KDTi//lkk
TkaGwoZg+dwLx8GVyPPxrmCoqHBHXwfXOBVi3f+V1C07QjM9mqg+Sxn5UkAPhstl
ki+yf1mVZ/d4vcUzslyt0q7WLw+PsF2YwoI6NokfiStL9xX7SlT+DRcqaKGft60s
dRy0iTE2IB2UxJ2u79M+yLLmjdJzbc0CUJz1OcsrW/DW0Ly3NhJVSWIiVsJKG6ep
aPYPgpVSx4H5n9Oio3K2ptOFN/xKBfJRd0gdJM9pc0xY5Ft+/+g/rxZxuYOXoM0S
SEvCXBO3U+GMdzGYWzdApU5cnvzbnV/Zo5dm8ConYegmekBipYJsg775QBj7B+tt
QXkfSJMVTHbJi//7jfR8CFe3elw0MrkD1ecu1F2bDJUVbYyhOIlptsWaONqN8h4/
5KgrnSzk8y1iC/jPqqgjkJDZp/BvjpCfRsQdGhRnVY67z5wWAhSPnSLcIFNvO0IJ
5NgJiD342MMI0Ul1NPkK+ro+FmcU8FyQIe+97yaxyVmIW6gDX/vcjMvsaM62ib10
v1ZvBbk3nZplpL9fLnQCLgXnxBAn21JfR8VBt79NXfHO6QhDvlGJOVThiov/ubGi
KBK/LLASn8jTsMjJSYJ6ygS1ohEQ0fPhR1udmJY+qjFxflIJeiIsd79crsfv8hsV
2g9wfAeJP7xgxAiLHlRKkz/5CAG74MKQda6sPaV2hW2RTIGBgZg5D2/3O2msaeDS
DDxBJVg/DSuJm+LF3vu6fV3xpvCd9eF142ucrR68oq9fvozXG2qoNanofR09UgXJ
aMwwBX+AC5M9AN/F7TZ9L7y8ieuJM+YopqQW/MTvTJt8+q2IIEdGAKTonmQ5NL27
2akQV/cG9heN8gwbt91d6udoFlwYGAZNrCUADwChL+qRR+7qalgJzPMKgU5dUUG3
HG2Xig+Z3f1yfxY8Wk+PwTs3Jimunw91MLXnmF2hAlcZwWpWShgSzxjIhsF5hrD2
5tdmbtiFimf4RkZVjxH9v778H1PNuP7SyMKyJD1jSHtg1ElCtyNPTU7J275q46z5
RMnPM4Yt+l5e4eCoq0WhZnoWSFIzABdqjAWT5LktS7eQpKaO+1up7sw7AiY27BWZ
95LUpqYdWPB7+cyCQPJKlP5ApA9+9RUlqzAx4OKwagcOcGnjc1B4HrRPjaI+MJ7o
iycOnNtD+jZPLZff5G83SI1t0ju/LoAnyb/208QZvcJL/FD5fF2ebfUpIfJmE4sQ
iauhkOx2YJvkOVTBF3e2ZXByxCokB8ivrvHol9YiVZryRiNPnKVSz02rpWb3swZu
sSP7PqJfOEsAbpUiuLvPEp30SKwUhJWXJ2Dq/wML/dy8fPcWea0LpwVDXDWPzesi
3xBZwrsw2Q5SFP5zVTK3/acALS8cjj3Xv1bEwfwPZ6n1w/7y1eKzq88q2W7DT3Ix
OCLtgkgcn2pvgAp2oRGqvLIYUnC+ELx/bfImL47JyvsK6Tj+flJ7BaJdaA+NwG3S
SB0LOB1VdjynDmYlpm3lTDVBELxd2cI0naduJZyrKr+QWaYZTpOKoRf8ah6c+2Ch
agshnwTbFONMjWSs6XPvHeljYOgN//oPq8oSPgQWNZ9pvQtrmRn9WiehEeW5zog/
iQ9prtq9J8Bw3FXK6AV5qCAqkM00NXGUZg6Spzx+Yuec9OhR2q/Z79MzJXlA3rBo
HazUkezfkKGNsPKxovqHeW/o0cXY8XGcaMcBytkQms3HBGz0UafL6DaBahIfjG+m
V9eT7p/GB2bhCae1n2AGv7vdxksmWoU6kYJq86RjjM13fe+0RnrNhD89uFyQSc7Y
7U1EXkp/PXuDG0SIHB5SfTUYtDUxwGVuwd4C4jWmyJmnYweN9qMh3qP7kBiuRCa8
M1FT1886u+Ubr8nWh1wbNys8IrclyEcOsn1iK+ClkiiRF45eau1/2b7+IfNd7wbG
+nGT5zvwOFwQMUqVZ/wY1+fhe1jHSX1bQC9tzRl+XAUwvmJIks7NiWFSdehnex6G
ZZExL1pYFKamr75il1h24UZWxHos3sMM/uBXPSPsQ236V6eNFi5B1QbyOFwKmK0L
p+k2UdEK4k1q+Wh2RboGyzPZwPFyrDcIUEeK7e5gLwVT7JaKerjDaCwww55PvW37
UZGz6f1tlovckNg5uwQdqSQ7taspwV3Nz6BZs8Yd/IUmaj+S985zBEw2/jwhZg9d
v64jDkuDiNniDd8dSWWHKopCYvjmHqn2Z+WnKH8xxC4SJrA9sPFmfgmiKFQU9Xcj
4tVHStAiCuuEin8twNHWrpNyRdOo5XEjPJeuGD/FmK593YTU9aa9NPaSYe4gg+kc
nV80mzanJjjIcxadOSpSfzVMTuRDP1Gs0leFR0MZ6Xnpwl6QdS6c91194TPzrLRl
byPRopS2vAiSExvUrKWiVmg1eByjAxSwrJwjfu3XgDDwZIsv3Xssw7lC6NGYznVB
IyzcTzVbQBQGnyY/+I2ku2S6qDdybcI27e9hSGUFC7WBqr7VWJcXrp5IbwsgfRQ6
u9d1IBNnzPaO15g7hh979r6Tz5+OA7IPOh5+nJPejn6IFDKOgdWrP0iYk8S4RWTD
5eYTmbdcrJgwmYxfYqVQDzYxc2ktzrSEhdabr1O4QhL2/S9Fug4Exe3hNtR3siep
APas84LL0sWPw2AOikwBroNFypr8QjQNxABqG/uNA0XDMkPI4R6OXOSldDwNPsbi
Hf5XRMjGz+TLf8hS/58ztSB0B84lmXPNJMgJiTJeubtjc9wdQv/E5WDJVPIgD68k
pVhdlxzCTp82G98/OPgkst2tTLt6nUwgstippgT7DL7OpV6l+KvTaZTf45piPWlU
nIP9OH8QOizns7RXAfFPLSF3DJrP3MQP9hB/PDVFSgWiY9KhFy+35tIcsxBi8Ahu
jjx3zwHojv4pUFFoin03oDnMKFCkKfdBQwCyJ2yYm0aI2MjNlgeST2hc+2NNqABg
oiwo3vPoaPVEqeU9h2o8rFRtd+LflI7pXZHbWo6kyBZ9/cVOVUQIi8DSHNOAhfun
Iocc1IXNk7qKVNokvN3g3VK/kqO8a808m9X6DbvFB0QOD9SDrmyRiMc6nkYlARyj
wYzh0YRlepfRcWf/bSE49IzZ4TRYj5lOkbPPIwmTkrkjenhl5zNCTWKdX6b0MmWi
BBExMUtzHAHAgGqXSqrdxSsbQlXI5WqpMRKyWy9HObVWHzYtpdOIFePVWnN3U742
hL5qjRGmNzT4XiUFNzsMXYI8D/FNtVkRYviDB8jTNELJDIGFvzirJi+6bBdbEvAG
oXkDIPossw6q0C8NvQMc+QNk3e32fvDe5pdCjMyY/ljfsB+G4/r1GpzK7QElCOzK
fslI9qVYdl9gcpUv+a+grxPvQPLB7RNhhTC+lNy3EU30xpnjkreLJ3GyEmRftW3E
j5VcyzhVVq6PW6q5FS6h3xikK3Kt5t+tECSJdcJJaLOQupbXFYSIZJbZg0k9Itbh
g3UG/kHQ6lutUmLU8C4ZxopFmpikY+bH4PFMzsE30ObJoSTio3GC3gweu400hZhL
j/ihyE1MFXTGUOJIaT4a3a2CuWmaekCIiNT65THzBNWJzsOkWAcF9Oxxj5UJwEyb
DUjchcGILWRTLW4+qZjKTh3aho3iLOQLtnC70Dpoa+wUyUZOcy+7iM0Y04OKYQNp
dRXc2C1Ns9ys1tKfNcqpFjs4aO8ttxT7nGsAlXk1X+SKqr+SR0q0I6eu9dJW4CBo
e/7YG2bk3BbCGNfnuWvvo8ISPr3Hqyznt/gB/BeAiT53WoepQ16FMIK+Zoh1YMGp
J/ymDHBNT2Br0L5pjPn5unq4wNKcma19RQ6vZVuaz7lp1KxPHUJVxIMZNfv0GmDo
nOLQyme0J/XusYqkR+szyg8+Mk44whl8Q3QewHwaOyld5PEYkpufzRVix65nZMrN
5/OowNVKcIgDy2KtVR7ep4CibObBsNKxEDEIwzcLU2s1lwwCWOAudObsjUXd19DP
rBFqfaz/mKcBxjYYyTuVuvQ5RD/AWZu7EDhn4//RGDxfi6DMQZkVyRr6dF5coB/2
qBm9dXHLGPrW92zYn2AhurXdSd0L3rDQfjUGr2z7EoxTGHeBTlwUJj02DYMIwkxX
+L2DnqVUwEaXNjxiYrOAjkG5jkceYH9tlbNuc1J8K+NN7RbjYY9vj1glu10ak6aK
kDHyzh711rOlLXgO1PwYINjGawOw4944z3Dv6qBMitNT5cK/bd7N6fa9MreQA1pM
ayFZYNzYxLHBY/9Kvqfbjz3oe/M8RMzJjLBxgBjxeeI3X6cCS2f3tCZoNKC8NqAM
IYRcmnfvnsG8+iZWVHVkf2YMzfVjSZUYGSzHOi8eFwcFMR6dQ3Fmh+MPWCn40nTu
8Z4u4NXu3fqOq9l3mf4CradfSANop2mpV0QwcW1NdS0X48K2QH2ryErxIVGZ3Mvc
VXRkBT/UqGHurhGrYl5I2vf7f95xK6MmIM8R/J5xLu0Q5EAqkGGYN58RsVuY0A+/
JOEQhKKg+cpgHnDTw8pxLZusqiRg0Aw1bh+7g/lkhNQEwaI9e8WTZ7cP3nF8r7iq
mPqhlEwwBwas7juYgx4U+brIK/1iF313UK7UzoDmfcFzFh2DBTK0qmSU1cPdpdJq
9h3eJ/cx24j8QGrveYYiOJvhFOSWYiKSINBqMjchXZ8UcsoiioLeRriVtJApq50d
ZvfAO+ZQMuaHqXgH4nKWb0rl/Mm64gi4hAnCP1wQEVmg99upaKISW9JtwYF6O7ty
nNaf8iMD8EBURsIAAQiHQQ8h9R2AghGKfljBTXhU31ZrKzOs4FghbQ8D5Kk29DU4
LoVLocBQp6L6fwhsi1VswrgjGkoKzv6FpKgfDVE948qOF3GcCaoR8VLrj2ESq57v
bOS0wyL62tFJfhHq4/LoUerGUjMsRwvo25Is9jDwHKCKbXLPb1KnBLK8gNZPSyTx
gBPX5+WBlpkjKYXwfJUfPRPTAVg3lA5A/7yaGeffwhESBHduevzIPu1jsfQjUBkz
Vfi33cJdKUNaNo8tPOgGN/jjQBG8IorgGNHk4Npc4+sujQ1QZ/j2U90B4DRNlzoT
TeccSpjq3vCL0MQwbhCv8z6QFe0mU2WgrqxnxdN5k0eg85505/Rki9453g8DcmI0
/fcmzrx3yDStAYGKL99Ur2PhkVjgJ9MASRbPGrGb0C/LXR/r59Jb/n6KVSoor8w2
cZHXmCIPP3i+024+hC5bweIAbt0ATEoHSkSh7paRBPAcwrNye/T8P717XIauc/0l
x7g7Gpk75/bWEk0eY1czylgbQpHl5WhBDQFAkpLnmp3kiZ1pQLwwsJ0gko2Z2aGn
UazIeEMIhYveQtFydLDZv8rVbMUUxE1cGx4XEtXbQR2xWF4cWuy6d7YXZK4Du+NE
gQ0VeUBX5UjVbgD9JHqxX3Ut5iiXrj7CgAwBWJGsva2G/NPBLWoT61WkVsH2VWrr
AoM9iJbZ1abO6b7Dyi8F/4k+RbyNsUjHsPAkl9UFMsoXzfvZeK9jq1ESI2vrvLfR
cF/w1j4KyQFq88+g7uC7XedCWJZBuU0P2Ta660FdiVahBLpvDco5Y48rb7cVhJl+
l5tMYD5/6McHB/oxkEJamL1pdmMzllimka6pPmOuruXfxT812s/CCa1PaeUoNlhR
RRHrmYDKdBVF+ie2G3d+64VCbAWKQathxMKo8N3cFLD3RJaEOGDdfcjbb9zBbGYX
x9EqKD7opK07abDXMZ/XcwskUxYe8l9oHMqwoPfR4wvdTximICK89rKnLRujnkHE
TeSgyt8D+Bwll6KK8GaZ27C+DLRYm3J9dOzKkNZ4dwRpXBX01+4lQ0QNSlaBwiav
Ad6g4eBd+KIAS4NwMVMHBYpTHBFop+agSKh5C6YAb1xlVC2LoZAIY5ucLmLaRV6+
bSPPQHLpdXnlHbj+O9b4KwWCK8f3OUA070u9sYfDIDmG6JmFCrgBlyVsN2BcWuLs
SzFSmAbF8//F5av3ax0Z7RA4v1P8XOqt8oljlu7jCO5LP9+SZvXGZfPnLEUlDYi2
Y/nzpxQ8wNWP4m5wNGTeTCZgMsMOBSd9Ot3MOUIyFApIDwZRKk5xp+exqb+GU0ZI
j+RyJwJA4vi3dxgAcpTADXwAmcCIsa0RGajm2PuQ+65OsIxPMi8p/x0m9eW3C+Es
squ4ObAzYWUjnIvqHcDIpISaztW5kY0Fc6bolVPO+nmZ5nj2764XIyHM43bQshX9
sfxE3SGNSY3YmJQf7GoYn1lPQX1PlxN4eMmmTBvnMhvnq4KYDUqv0OqsMmvpWJ5/
lvOA/nG6JyVvfPqJO0I65h81gYl7y45BOIIhJK/L4dojN6r77N8ki7MGQpqF8NLG
/y+QcISeBiEnM3tBb8fXZM/pW6zMDonuoKoDwawe0G2WtGLVYAj0SGjTnilCBeYw
StCRrUdJZBjquHAvlWEzbRg0Reju8EwAdj/eJFCj+aRntGQ1vAD3dmpG419hR4J2
/Y5Za1YwcqFqgf6K0+npZuOZBpj+KP4/ewog0WEZK6B54On0gCzVah/78AidjW9j
MIZ/6fxuh0R+p4VRGCNQFFkSTuJhLg19N04jMGnl567/WykEDwvVrVFduEM/CbyM
vf/QslSVtRejw74Do1eSW08Ml6iEogdyGEbt3WDmsPVcxdlL4UiqB5vbsJ+x1JFg
EQbXdZAwq/tnCL85RrNG6owXG7ZZzZdf3sZWVX07iN8eXPP+qVibol1KEhJC4k8g
GFJnVXVaCgOkNSoJ5LLIj9qNWmsxLaY3R5IxuwNgwBkbyl0ai47W/K6lYVyKYYim
Q8RgT9441qeGIJgf8Fc81gMNCPxsTALD0gdJ+c6mBBkBRGwRAGU04MHm6Nj2sczE
6CAn9CJPXoDNN1DXfkmL4/Rfpc63425jeh6Ddi7cAZnpnQtXHi5ljxS0+2Rb9Mby
OwlnTYKA3lETNM+r2gDTsW8776JFTYL7/uyTDEBR5HSKT6LhvQIZSJ2to+u6HhcJ
ykX5b7WSwFrr0WULFjf+ykQN0IfKoj3VRdqKdHSUEF/q4sJJXsb5oYV9s950s+La
5AmGybb+Qig4k7P3k+p3E0C3+3+TD0sS0eKqjfTsqNIwlTPXd0HxKV+fqcvQ1jab
D4WX7VapbIxtJeB1vnkRgplII+gLYYK4nmwOP8V7yJuk3DvonPuyhUpJvFXYevu/
IRnGCww9zw7sHXaQOJMsZ//jShrPlGhq59q1XfQ2Q1dMYbM2GF0Pnv3fjTfDiyJP
La8iOzFZ7TpwNdl556xWsGY/kSRyBQh17Qm87ngddNwW5fxiKV4xsTCIYsjfO3XB
SyHrOun1qzS0PdXAED6n7JrxsebL6SZUoVqePRC0gLF5Imx3/Rr2md4JlYJFco0G
8ut20838MX7+Jc+HBhrPqd5uPQ2Tt/psClxOXPogWIqkLGvBM1FeDqCS+h3I4kgj
r9nrt5VsctT/YI1fHNt1woavJ7JyVnqaqcGYyJCAIpfiiY2cq9FrdoTteDyJn7mS
EtJhtxAdpIYMJYaHZmR9mWBRW6uM12cXLoIE7Oo3P50Mg/le2Y4DkGuVwmYlQxcx
opTvW/DZYo79rjXCXuMfg5IgdUxe5H/zYqauZIpPfkYocp7ukz4kND+ueuvQ4++A
grAgO2c8NY2g//fcHvD7WOar7o8MMibMa4p6+vkNxT6V7vU9H7gK54j70f9gjL9j
Dt0ygqijD48BhCtzDop7G8oyIsDwyRk/SqneelcNcpXu11NC1QjjfP82WLY1AuVo
f7jDyQBs9pLRVLQITZRqTrSJZB84qbVLbc+OVZwMbJ1Ryw3Way+eD5wFTfr6SweT
SVZAzI5ZK/627dMjBZ+I7p8Ij1xxVVvU3/vJCOwZt3CGT1yeIyP5XWgeuPozIiQR
Mzj0gbprpIqHO4lgL5xMXAxGnwCqOhjFTKIMAerPB3HxdBVRrptdXwC1wT+Fai7D
xBxB8MQOx2HS6eiAIDt4IkffOu1rRGYY4c/uM5dseRYgGL0xkeOBPoqsA01VlnmX
KYQ4gEWv84yrsjZ2iwkZYClpFJjbK7RShLBuxZSV/ZRIOZrqKC8Gc7WHDmp0wz3V
IuBLw91Yv4kNtswSDuWvV2ZnUb112vi7K8ICdH9wZaVpZP6WdH0ZcQO3bMghx+1c
CDC8OMsG8XIB7WP1QNwh1OyG9UsOWcHY8l+5fux+HZS/YXp66B1+IIph71ELbK/o
kq6LJBsWzHFiNXGUQGwIIC3oW6L7TYN6zwyFzVZgHRN+DcIAeVdEbKdxoEj32EHw
PYKLv6gKG+gkY9ZgE4OoeGzyA42CxQsq2DjO9+FiOyXWJgU14ggui7FVGn0IUG8p
Kar4YKmQ9s4MdHtAeImo8Qb6MWVoXyg6BCAk+oJvVBm/kyGWhrtJRiEHkYtD0ATp
+o+oubIo91aG3SAeXF5ShEk66hUeXD8EmjRcG/zxKkedoEBa1mtEuob57/IRZlJ4
4oOiuLHMIuO+clPgR9XLg9B2EC8Q5FOjRm8ATEux5X9Mvw7ndmQb2ykRkfYdXgq4
i95xXwfAFVQIVE81172C6OyIiurlp8mPrGxut523CuMiCV+tOyasqwpfeNiWuVDM
MU8QqNmzl+Cnbo8N1F9k7ItmHh6WkM3LBkL+zRr+xxvgDxu9D2nzqR5V38OclJN2
L3+ju8QHNQCdPtG3hme/VLpjFZp84Uk3WAu2nyDoB9xH6f+uJuPug/8Wp/5eSu0t
bVAv7CM2+f2fTfPDK+wvAID/JVqZKGuvvUztY5bY9fkFeqfsTrijnKfGqSKwwy9j
uFJ/Hk3+BFRJ3BMFeACO3s2JFKvXaZy+CeG6NejsDLRff8OsKeDUMPa+mtH3WsTa
HaEVkbHrHxYTUAKkRwA+8HHBrQ/cv84DqISPT3pdDf5+DVHvJDx8hzqxggIgPySq
F4QKQtZm1GQHyfJjPJkhikvSUp36dsbc8eu43Oj6t7csbusExhP9iZ494bVmKOXd
y0YCkGJyIHcn/YZA0btTBjTVUoJcFyrZ2uvBxfV1aaZf8i0PU0f0kERbAW7U4Kn6
SZRdyrkpGjIfoCXQ10mek6l9AWqG5yD0TIJOIS9b+10Hj1c3FDTMQmiBkHGETI7q
GSL7sWviamoLQCQ72DemoXP+jgI+hwiTvcBglbdyp1pU8IyYBYNOdCcnnFJGIxlZ
3eur569VqLjDttTZtWxQKnu9womyF5uy7N9aUGrYjJfI5m36VEgyzj/LDFeC7TM6
C4tsUCgATnc5T4D1l8U0omWMPiEH/x6WiGSgBFssSUZY6K0VCvAkjn27KUrdlG7d
4P9Be0rIxzSHGrE+te1JqtRTz9ZYWznE+0WHkihBz6IPTB5lFF2RjHtc8INIMqKr
UFqcYUUm2ivqoWD/wkJx+t3YX/zb1quDjFQDztwh9z5fVBgTsvXoop7mc4PoObx0
pfPvDvLHZFLPK82Y5n9TwSY5LueBjnbgN/FKjOGAycJP2NN+MTpt6dAozVAZrgUH
Gj2sRHZRf3t26o+ecPeeXqeYZrqt+YgNA+ERkqq3hv8CE3Nz1X3ZvigJ7b8DF16l
LqbjeO6j2fraV2ii0NHkRWcTY3iEsADM4K728PqRgF6kK1ipgA3goI8GjJgz9jbu
TI/DkuadBN009tTvVmY+sS0YcRxds/FGNyOOeFS2upgJV7LwJoOhmAIrHYkQ5TeX
jynbfLGt/PnNjfEl9TxZlw8nUgRksrxSdIRiDAtF2DgUPV+SHbBMK9ZjQHQF7qdg
btDXaw2DOrixzPPBbTC3pIumwse1z6SSkxLOQzPpPCxZ7KjWCCauEUkrSjcQbi/N
bz1/BnRi/ewORYLw22P77lXH+gM4lrqmRmRvwHHaMXEZcKo5HVMFk47aWkMfI2Ay
yJzsfeJNGA3bN6LpeGTFFYiRY8aiv2y56H0fkgnWFI/n62x3GYdYR2Vgf1HRtfAq
5ZVZIOa6NpXFu7kSKBU0wp7kYdvRyiMmI5lw/pq2kWuGGRUFVHuRciwOVfFFqBGe
DEAzjjErZFgykL8biX87iyEuf3J5GEXSphjH6taIgFQvSkPxY5yrFaZdb0aQL6M0
zUtDPN5msVxkQI0d8uiXOXLel9OXoxqwkD81ej7LSvoEWuCwqnvm53Wvcrwnz7Gx
U+NgTt65bHY/tbSGIIcYFGU9raFXwo1ewdwWlbwIUBnDAxxYxmKa+WHcCjHXLosz
/w2LWnN09iRfjkueJEwPYLnBBazFipnnYM/qdNcEjCx+Y5YyzHR86QAoq/T1zn4V
zO1tuYcB+AzBA8dFtcgGXTGDNRFZ0IpFVkWxcxCyvKTwHxvM8oxTS01Zc1XMpjVe
ijwsLKnqcmcVzxXa4Cc7kA9m9CzoQ1XOTHBZVGvv5UREEwPbGzD3GuSjveQP5YUp
sjEFQC69xjnsIm7dcBk9f6YmCAYyJKhwPl5UW72gFDHsnPUiMcgmzNHkx0bzyHkd
1c0nDdoMVVwkVn4F1N/ZIxnQXPk+i+uLKzCAf+1Nb8rvYPJuhTJlKmMXogOrUqAV
OR72FYL6KvyE8hqEs45hMyVmbr0yB24Pp19k89lw8327GhyazkUfhE3LfJpSG2D4
+zEp1C/fAUDGms5cd9DtMjiLuLkhJcBM2Pk+N4rWR9OB2/ujTo2+ppqoMfxMotyh
0jyjDfEYc9lTgE/d4iTA+lofXCG6IEHp+HSnbuVHS0VAP6L/EWtsD10pg4ZLHUxI
HD3NltPlRnTq9jRMiJpicflLplyBmJjmOJ1YOJJsmqOLE+Ff6TzxxbBOSYmEntC7
gR/CPLtDSzNf7vO6hdcvr1gwafEM/aBDaHXLt5i3L9XD8MgDjOCUX66DBkQs0I7s
S8W/F3V88rf2WXnXB/tYewWfrFxLERoBTj/wCX2hRj29+ordzhrLg83lYXyQpcHM
N8Odx6Od1eb9vl25cQRMxCzjpn96+vp55beHyaK0CpQqaVeiSzkdPJH1vH6CtTx+
BYKF3fIm8lTza84hNLK8hrnmuO6p/vyQ5dtzZJLganOtKPoubc1ifDL/5BzAzRxj
HiDt94B1Rz3KXavp3Q3goh1TXhSunri4klP0LmHIagaLYWKRNUs0xN8fpF8a3ECk
VIPQXlfIJelH7O4lhQU+OtI9VwL+ZiEF+BuXjp55EYdJxvJQfePgWEHmtvIXqKJi
lJqT2qz7jZD95vysPFbQ3SGFJpYdPoRVXgzeCjsLop+nAWMCzNTXraqU3tymB0LU
F7DAitYQUs4JiHISogcXWkeVy/gfQ2R8E5zQ6vXxV02blsW2EjhGCvcVDIGqvMQi
eE6rRw/2xttmKGhg3K2XEYLQd7y/4iAytvg94hSwy6OyX4bPeF83e1u7yohm8KdR
zQ05gJxBzlQ1ThWfCw5HsL54MahqrjC7E9zGw5nUsgs2u4rhbwHttSP1xOeyDX73
RXR7c5IlQU5l4eO9kXqk/6W2eVEMrYWdS9LCfkRrKUF0ldU975CNYvsVx4Unmz0U
mzI4ZhllG02I9SIpz5v/XqaQtVDdjpmf2/rMLfgnqikoXoeAgxKZQeVC3u1LqeZI
Nnab6IlX5Bm2ksFv+wwXEaIIREzLldm1QKaC+kceOyU6XAAoo7plZPAROLuXikxf
6ncwDCXGYmE86hpG7JaIFOHu57+q1wfYNlvS7cAwICJWFAMOsrPLIGdg2cMnMIk3
BUkCtm1RQOJDUBgpzyiRxJdgOke+RI6Db9mv4LRLufAcnxddpgIO+3yGcfhATqb5
GCb/NHV2srKC3fQqmuj4aM+zfdcbLW1s/DUDfTC+ItB16JpwkKVtpm+pnOcJ3DDK
kVAzs+9EEYFkscvDFv8dRF1hBmDfyAcMWSA7vY5X3PszgRfuauwQ2Z7yjj29UAD2
xnKLS1UAKrUfWBaInJfR0/4KhwuOzhLUBAbynnjdldHU9aZGS/Lal1SkFG6b4qYV
zqEkwbjQhvWO2clo/oalAMVjGbI2iSrtQ+1F+8GcxXp1+DvnHRxCoGOa7erOMfNs
9CJgA6YVSp7WFwaSkCYSlMhNfDjQ5e6YQAjBG7qqlkQGssUmPs1xUlSfRVa0hBRi
BccYm5Ptl8zdJBrx/Tlrpu3VQWO6sAuBJDgEdY5ODZYuIyEDcpnpWN1xbiE0/7p9
SMpYxGUmsXPn+c7S1isVPNHvg3zz8nCPu1Kv38NKo1sd5znC2AKGc8bi2B+sIr0s
kjD52qOiMSyt+kX5VY1xLOVI1tsI4d+EoA2wAUQ+Syl8SLY+FSoX5t2nS1KUcWHn
jKAlPTqeAz7haCnwy6Xb3irZ37OBVXFIIeMFgNihuKKR4IkXiRHqis+wDZbX9o3D
yGp/eCi9k3K0NwmNmaLjSGBfWzoYsU+76K4T1jB5oSE5oYsc6bGG7qLT+UrOAROI
jA0yicBTfHCMIGgwDlwd1BpDd6tcSCvKVrQPVW23Kon5HG6dGV5PWcH0wUoZSbiI
AHTvtoS1BR60AMa/98HpBmR8xar6bIzfeybu56LXmTwlKq1nC2NlXX7IbDtxtXY+
tU7rYh7LT3/tmdi+u7rq9zhN/e+DQ6IzrOT3vOp9kaX76qA3VS6oRt2vKagaVduL
c6xScie0CkekTZ66xovrJza3Og38c4WMaOXBPZgi/25Evge2xA36YLkM49jl/iuq
TDJl21Zv1cqN0iHM9y0TMAOYH7p9/YhiXCMxkKW/mdbIsAtYMLG1iehmlujLbgw6
zDntLaeBCChwsNTMS95U7c4PwcyQYGTP2EeZRJKSLj1p2YabnilAruIuooQbaN2i
cOxF9HjJyYvvDFFoeWQDyUROosH7XCCvxeIrCAy/5eH3aiNVFcMHMdnCGMiBQdRp
sqM1sb0A5aMTLL5qz+19XSL99S8qRlZjL9NM1m0DNVmaHulrcMdhYaYNC8c8kLuT
RDrjkoAsZf095kZUm15qMgBqBFCkmUlhpnY3qF4t62EjuB9qAV/8JXmDhK9VlxQQ
tgg3ZH/Ppd8ygJeQT0EJbKjdo1/xmpSjs10kht8PTKpVj2YhQusjOPD1NOze1oWG
vjUn3sXKbfji6mRruIOENkZdWx7id1s1nX35wHH+tyt/py+DFuLgcCBbI3bhYwhI
rhewP2lEkgsO9CCgZcsofpm4ioj0YNvLT78kZwAlLZjYFscEFTYkr07o1EJ4yV8G
ri0Wu9MZzsuJpCzCu8ameznQzeeCoGFMIBUaYxXR9q+jaIcdRuBAyUgjt2zPOw2j
E+cLxnjQuWNSCtidcJWRcAoZfLINMdLnBiUYhNQw6EwtZCz3yJIWYxSXDI3dsopu
upFzt6XY1/LMkVkmKezGRDjs3nXEwqqaOeb09E9vx1j85c8ac9KJP8eQwHoQE+8i
iAea1FuPwJOVptddfyU2nf9rjDqsIiw9uM20BRP/cJ1/cdpHpuMNQ76u+/Ej4uau
JbXz3fGXe1tHr9LZgJM6r4lcsLvoh0CfreEjNIF0V4+1Eo7C86h5rJGJ4AvqM9Ha
O43LgW11KtHL8OuSMmLrELWPopWrzRTon4DC0rS9MBpk2vCn9OBGdzk1K/yhVi1S
iy+0MxgIi4GZzNDA35Jr3czLawkUglzTPYsTbUCR+y6L0g6BDSF/XiNOXZA71CjF
5NlTvZzAO7QlK7XWdXalook1TjeMoLs/u/40wTFVU6pS+yAAPA9ztQrjh9BbvHSK
yu/O6peKjrKrANIWtk1mtePpkARGJE2SqRgGy6rH9BaUD25zF89xPnC+TPuc0wjy
onphhZuid4XIRKO6pJDmyqatGb4O/q4NpW90F1OnLTPeiPIeVeNfKMdERB6xbGOb
P+gOeGeiliY+SiBr07zzPLhv/cHtPmftHQm7Sk9Nao2HXoSYXAdX/qOqshCp/5v/
tdtV2GyEU7g7qSi+pzEX3mFeUxzQ2/7WXkemWU8lcnAE+JRvD33C9hzKXBDFreEM
oX8Gm5PmjXKmuHINMl0QozS+u1XU2iuytabr3EKpCI+prudc9pL92uRiKaYlINdw
PI1Qc03eFdSbhcDotKHyvGJT6gogTPQSvB72DsJ5wl4RXHFWxPNsSfJJEwtx/QbT
cAWHH7+jGLmHxcrsHOxqKe47lM19mrnZfWzM45s0rQFYE+ClCgjdIsYxElm4+IOG
Qz7Npe51fnZ6/MURtgAW/mXtoIJJXp5wJzorhQ0liS8/oYNqzMqQNdXRC5BXXRSS
4MewilUT+It0Jro6VJGBSNjXlkttTegcn5gCmC6jIYpV81hAuWgn0BvZg3/9J8ta
+NuWT+MOzUJ5Q1GNPnw9MV4IG+mUbLCjBNLeoGQ7/bYjK9LYeY8vascxu/VFbi8f
I4cWijMQ36mKfnsoJz3yu/0MBmoBcGSO144KfyHKhNtBSU4c1GsCH6H9h3AxKgsN
uomFBVOOV6nNpFLxLEtY4aYc2DgfHnYWHR330/c9K+In2JQKuUNU3vALUMmPg6Bc
hDqXKK5H65Bo34hxrRotmblPs6T4A884IA6c8Dv6cl8lL3kvS6XPc/K4i1+L5yQ3
Z/zILlPcjWyy62RW/P7g2ZMRXhaXn45uMxJloIKtLoapsaF9ew0Ru6iIeLhr4/uo
jsUmNKXWqCVUjRe6sodWOq2LMLxOupVl0+X08VBfy0HjXdPLbN9uoQF0cSC531j3
bt+u6z6yyVLZRnrfl+Dq3NeHIIYqZSH9ovB+j32iqiYNaD4gpYlVFov+M/KSSKY/
QlbsZAeUVm+rD00QMQgCcncfl7nYFQT2kDPIzT9c57p+2RoLG9f17ffrbsP+kOp3
ArIMsBKC5x7/qX/Z6Ed7S9OzeK8N6K1f1QcbNxR5e8oPw2N/8uwhMXbVp+G0I3aT
Pp/R86hvXBDUmVUkRSpQAmdloFNNsYyZo5D6ALM/rvntm0Gre8kRlJTLm3pdFblj
CAEmmPIBilDwMgYxxYvby6tb+9utT0Bfy+Ic3Y1jR7fdT3mE7FXAJlNsFsy1Y0pq
Bvh3KviyfBTmAXMMMkiKrNQjpyLZWJqLK+Bb0w5xnQ4Lu/8M42wrpgpmWNIEYgac
5Y+bao3bmEj2bWZVGuY3tD5PLnR/So7W9UjtbIAW3T8zmCZmaiVgaReUDsgWU3rx
LiGz/mtTX/tIDmOHFHWULJOqCGUsEMCDueCV3Ja5mGwEvXNRUyZ5zvYYeEiJrPY9
hz5LNCi3IbAEit2zmi7Uq7JRJ1+oK/6HLuYX3/ni4NBkckAu5lun5/WwXI+5n55e
mrEiICG7JGgjkpCJFkbG+NYWxfOIVrq2AiGy27xAft493LZ3Ww0M7lpg4WDGNc9k
TjgmloBBxWcxekBtAWu1C+qy/6uIfrsGTbnI5lWZvbC0xdPpwnywns8OgknoADo3
FU+aFrpjcdVLBTkE7qEjqWm+7c0oa34hzVtpwvfW6YJ6+cV5WqlXE+YNYoWzmIrB
yTj6QN6YSZiXMxGnyxrXYClNOI5jH/dLeFSLzeEZyRzf/wJG3eDWS0JuY7Dx5aFK
k0DDffj45KtSqaQeIgrOhoXL44UmGtvcQhU1jD1KUFAUseE6KI2P0ZyTFvY4Xmde
wm1ZKX9WkKfJHBhqrqleB+nQxed8B78VGiHRzBxzOSRQTm0DhE+FkLrrYbpvPp9d
vHLsnhDzsIeRSH0HkR5gBB5pNVn5jLjVMrLPGvpi6df1P6f1UZQ2jtg+vs7gAjix
MDHb64vzN9Qo5lDLkSldyM8gWcait8ulBdpNQN5K1xrYV1sVcIJnd9P0+0a9aGqz
2usz9FC6QVlL+bc/YmcEE03AbYMnqkl4TwoMB3mBq7QdVsJge5q51M0TCNzZa9b7
ruq/1B6OvW9eE98t2ld3DWbFnhOpju7Gzh95J2lBk3f1f9OhrTXMI1LtI4OQq2wM
lWT3lcI2OogLU2oM0bsU9FAUm+1LLtqHL9bpwwuIWDb4yq6+pYakQwnq5zpr7vK6
3SX/R1YSaGkLDf5+jdv0JS9Sxb96/AZw5KGlSrwE9bws7WgeeIMUB4h3H9uZAi9I
gDHmJzRV/GUeh4pc66uNN6I/AzxvWeaoMKkocRiEglRuzCFSZIIe4ldtlZ7go53d
VeZMZ4Ta1/lNH7AsOEX18oJfV0QVbV7/xzyKO5yjUx6AhI/8vR/4LxbnRtA88isq
UqhWveGsv8W2wrzcoXnB2lInqgAQ/mjOmKWmxe9xFJ8dZCxf+petpJbFogIB/VYP
IfZc7oo9ZLgmXxWnNjngkp7FtQu/7Mp+oRgvDTV27P0INgMQpXVnWoniJy/6ecW6
HVVNPpgWYOQCulzCX4vYHSAQ46Xqv1l0+T+k/FPJ5yC5LiF5+/zmwDJhV1KMp399
p72vMEUJ/MACMuBnXAEFZ8GOVzBtsgMHNdaFeXD+mqKo9Zv1azlP5+R0UhUWVClq
TgQDsB+IaNziVT3Y7A6YA7pIsqOdbVm532Rr4WKdHl9y5qE9tEu5ix+AnVIF9iFL
Ckt07D+Ld+2dqTiAmi9WsP3Y8tP0VxUW5l25W1f94El5jurI4f/OeBwc80eDsGh8
OZJzC8EnXMjCMWKqKF1Bqjw+jtY7aONfjbCSkcNo3DjtQOfQQwjnFY793Vg3bylD
yMd8yqZt5SJMUBmGuWmAVxqQRJxYNP8bhZdeGIn7DiDi5FlmePK8Px3ZuWvu4rND
yOOlfw8apiL+eU4bOD+SRT76P/evfV27m9wIMJtz5c4RbEIs14E3O/LyzkQ9G8dS
nYDbmJS9ZGWkj2j+TSqCtCmPbMIkU9JC3IGDDfBCR6aObmDI2hws8iHYukbnAn4A
AKc3sFBBjfPDRmHs6rIjbz0k0RDu3uU983B6X3DRcdJAuWBctOpl1l63aVxFszue
Ztl8yWpDbzdHc4YQRM9VKm3dA1QA+kTPDLQKYFCp1QSWgGGHkrBhZ1Se7oKNRa8Y
HaDAwwUfoF6ibKHZLMLPKAnnbIfcpAPoV1rBrAEdnnuW+iegk1HLfL5KbtmfolMJ
b/rfVoYG/P5rWwdpMvbsRd2GRzORvHwRO+IGbqDEsM3QwUiKqwFQ8a793LdhjDNP
/UAZ1bte5OoEF97KTSbg0UcwaRNGavlz047xj3HYZldZUX6pJWPhjW3Gln7SbXgB
PKzcV02cKCXpTciWeZgBvLYGTfHbuhXCq9Xe2o4z+/bj1lGkx+UD608aBIZnWL8a
8gbzVUNVxCYi6RPh4Qa1e98zuT21fdYWG02vxfcpVxCke/q47Zq7FXj67/EFsbUd
jzBAw6DO+xmrvsnDZlQ1BYok04dBtz1amQem0xcfMC08QuTls3159+q+8CNAINXB
GudXHBTLPSEvoCkXRgm2i4Bj1YEEqqP1I0ChvQeF5zo7uINbRgrqkxw6XzLz6uCi
xuKLJRM6GGYbCt0ryOlkgmVyJ1APpRluqYxpt77CJ0zjnL9gyZrHXegEBqsv3aV7
QkgYd9JBS2z18sbLDmpiLedU9vzq7bUeoDxgo70ikOZc9QqYIKU4mjiOF2AR6ZWS
bwZNP+za2SYLRtMvuA6NjDmhU/zqIcw4VaG3PjD8FnbtyMJVtdrnKm8QferKHfdn
7JrJpUbp59gsSAoexCVpWfBdrs6hS/NgFnof8zlhnOOTZ+EVAtkwCuf6c3ICCVMq
bmL8t0mDXioa9CeljVAo8N1aaUwjdM7KPQ/kgtKTaLFxM6wwJfI/BGU7npAf/jxD
9NZT9CGYLWCdbYIoziXpueVPGlQYk/rTPLHW5eM27bjaj2m6yYaPsC+UDcvbQN8K
BY8QAVy2I+taAHPbOQx1/j+Jrl5p/RmUbnpXLLqWiIx3nfBKkVjPAYS9sXTxd0mg
ky+ES6j9oOYRUh2OhfTkCDLyro1P40f8JdrcckEdp9KH8VG24ukw1A2yd6xZqlGq
nM8ThmXyYRCtbDBOL3xIdqzVF42fG2P42tngYL97B8hdAsb5Qr2b0rj7EC5Z9KZQ
h3F0vYw3+muPBm2U0evxsS991GnevAVrmOkLvXHGnVgJHpQmS1skbZ7VMVw+oE2w
ST+5QM+U2ge9AQnOe8ppr1LiybRQDOc2FaCo+xqW/QypPriQolDwkdwT4R4BQbUe
xDGR1vXmV+nSlyMLld4FXmqBUiPNJgOL0bGtsUm5XLKeo1HFsdRXFrXdQatj7wH+
hJKfrUYtH6IaT3pRj+Xumbf/U9o+rGjg58rhX796WMKzarghNilAAycr22xYpRIV
4gEBdKDeELRbde4TwoIi4iM6FXO7Pb7Pyht5NNkdIsg8SKMF3cN3/JAeesqc4/7W
NdmdCye/SUx5Iv2bjyQ+ZFau07y1Jym5iqiNRu8AALzu8BQB459d5L5XtcY87AKq
/YE5LrELl2NTa+lfP1aEuo4XHEqJQg9+xQ1wIQoOcPJAoPU3+DtumhQpeIX5zUPu
WcfU+F8fWVbm9Vzinhcg4l8CPR/fMtBT1UEAP0hzJ72bh2OD+nvhBRidEIBh7VEi
PA4i3oSquVFqi4t6QMQWEDLauqzQdqsr+XbkTv4WLD9RCoQdKXG1DEQNiVpRtzGd
4OCF5jXQUEcw5HlJR88oMUMF3Ojo4L8wSd74HXfglaONAs38rIpYSf/v/Ud6khoI
EINCeJr+jzXjZP+YFRlcd4W6cjsl/M7z/XhE24UQBWmvrmeoV/qjpNfo9vLdNP2A
8RQ2d2BsRq5BzjlG1ba/49ZLDvdh7auUVFQxbJGJrvuz4qXLzlSgDCpww4qiOiDn
HKbIm7QhCKRbQdTyHHrYDTDVIU3r7VERzSuFSQMbaBZEkrbi7SqZ+TMXXpUy1l5c
lV1hUtcK+S+WbfFwUdh79wbOovzKW31KS+Rf+TCVBPklPcJHg2IWkcd5mLcuXfk4
BJWTuQ4T57+7nRngt5jobqesukvyAIlvKbMYxnHBJ2ino6SgCtkaDBNwOeC8cd9R
vBsriLec/4FZXw/Tx6Omh2exNb4rsbsUEdICic3nK4Re7gUzmw8L+OhNo2gPaMoD
U+nGAqrBA/Isgjw18RQhkWyY6LVMR42u406YlJ5MoT3mgJ41WarNGBkVmrHoij2E
8Mhp1nGGZeG3HoMXDCydtjMGvl70ETr9mfjnU4tgE3HJZRalgQu88iGfOqMmL3CO
rCJ9duZgrqXlNyBWNopFQPidSOeUjjfzOMiGMwPsPA54tXHczHe665qE5wBiRjDF
OZJKFn4CXwOOnAU1UIoQ5Y9LtDyyz5NGMi+MIoGMx0RnEyZQSE+QMkR86O+ucWDI
XHSu+PI5S8e1M31EIovIKRL7Rs2TKjqtEaDPL+GivimcGB9hNFKN7JJJwvikEuVm
mRpmNN25wRc2frzam7vTvT51kem6QJaNHNiY8525dKwjVszXknl2QDpkqWWo9Ouc
zg8dfrFTIMzNOyy0DOfo+adusXnWinYi3ECeNZHR0+0YZG0et530jD3f0enFlYQ4
Yb4fatsuqe+vRulSavCyhPaZuLa/cAz9u6FNWfLrw3bo3BuJlEcOLCBUDtyqtHsB
WuMCbrSXe1IY9C/bpB/ljIKdbn79SS/P8SFCk9ax9xQrP8GqZ1WimnAdX7xoiEzk
gWwefmFqWnDSs/MZsiBnFqyZyCJO82dsW6/6E8iqaIq8rYVXPczyfSSoWrBG7ga9
TyAm08edT5O1QG+CrKd2jDAWvgAXU3P9QjLwJDXjEJg/f23KPqy36ni8wtVkX/fP
ms3dmSueb9HeCOmzwRIrZs0aBfQaFc+k9OfOpX02rlpMP7eHfx74qVoxWHTwnwiJ
nvj/hS9Mea6OH/Kdb9FP3LFfoQTukz4sDKl8hwswyRR1jY7uOiB+ubxHyYZptJjH
2FcudYe8mMYjEzWtUHomb+pnnTQ/NRfevngGDWM43Euqx/MSQrQpF7oLBp8ZNY5x
xkheJ5+dd88ZHZPZSiAa9qk0+p/4jirXZ3U5hIPqVI4HPhSCm/cyY2JgmRsyxd2b
mUAAA94xYwCQ0JZAjchoxqWikwRlIG00N8MAHo2a8+iUzmfbezznWrsV/oC7uESs
u7G2sXtt0P+LVoSEafmckuzlQnaK8Xtao5EEcnxIyX2wt/LnhJLBbhzmsr4kPc3Q
Z2VclNILkQ/33xL3DBB6F/oxS66s3FZoqpmd2cyCQdX+O1cZvpHWnppyUdNahKrE
toGXsDfnYy9bZro3mx7LUJFLIY0lj3ozilbKeOV4ieFZCz2blWS3I7mDRnrmE5Hp
lyZPKOxEodpTnZLIc4HJYuHZZzraYrdbGrTiQoKXKLwncN207spK8MT1Ah8NJtxg
KGXdzFFEzi6d7EzKLXkK2c5f0RNYCnej5gSfCRQ92DXBbiCSqbHGVA45Lpq29LT5
cQQ0huE85vyq/DVsaH1Ne3Watd+wTUR0ewtNI9x/y/aIbOopdlVrENGaO1Opzlkq
E7TcYWfb+h79pkEIAtKdBUEBOdMKmicfONhqYI1qZBjMqM4I/zMYX0xFzEWe4iqw
8DouDL4/DNAAAgr0ftR205cpUby4Ovgc9oCtuzjvRH4FesZb0vtZsk+RzgHkGQLW
KpwwyTlggfyu83pPlKbSggs4yCzn5Dd29xN12DPjBC+AegguFO9hHJSvSjyCttJM
B5Rrsixn7HYbFyhHozwPps4T374N0sST5K0QMz+UrUQSqy0mvjKznr9lR5SukYLI
5QBObx3h6oembfiGJSkp4j+5H4+6pyMpHXryYPUetKHmfFy3YLFgT+lZYt5CaSsj
mBVUNL/3b0RBjE6gyDzzvtuqxYgLyiLcaxkFdhFrOnn/+ydnXzoPQY0mla0oeWzq
nhASqf2wnUl/IGydbnUzCkghmsVMYdjXcGzjiu9k5mhBuga3NvUnmLrN0uWPRf9J
FuotA9Jd+Z90aRoHisCbQrZtB9YjjRrDrUrX2mlDjq07ZjcTrpTaanpYQqNH46yh
PleeLCyzriI+vTV/Z/3oAqiqIKULAg/7RGdWjq28A4hhKLXdUOU22YRRJs9k7xKR
bJcCiqoETXnk5MTApNCoRwUMbXC2KZyuSdmtn8/XspKwkFVNDQJtQleHZBWIhzsu
8gaCDyKgTeRmTaMIUCsroJTA9RyO+H0vCMX2klKAWzPK4DFfJaxMxbvkA87azJNE
phWINJamAmJulVJxJAYFE3PPhc0jCOIOLZFoO4IoGpyBEOgyWJV7K4tvHSrOnULY
h5LxmkVTk7dxKzBGCzuOLUzmQSb4hEDl9qLuh6dh31TieNlekaT6sCxMceSom/k3
e3msVZ8ggwKkrlix0o/UwEhV7o+k/g/wS3zBw1S/88cjn8UzA1VbFqkPWdLk5S1V
heY7aFrSHE9QEGhZsdswku0dzFJ/SD36WI4icVFWqMFK4f0z4h8xEp/PNZT8DFre
shv7cDa8rKc9oRxj/CcQrimmhSMl342k02e+8hfnYonp/NNsPW6QEmJsAGDA0D7Q
eUnSItOmBx28vf3VVB/1iAPL5djTmuowNsev7orchzBALxtZb+oo51LtAGScyIc7
tkwQ2Vsjr4qej9Nlz3Lsm/aglyjDm0Vo5BlTBdUygpVcrUDL4Y+jdEECc+8MFEAt
iFijkL9ngRTk/75rspc6CZnRuOqVFdOKNe+GYRt1jLUDqfQN0fQEzmP1nAo83wVI
QWFfBBpAFTwqIUwxHuC8NbgSj0Df1Wre8TSOKWHHVbY0C35IGv0MHPZbIOo9BsQs
WVdReTRrvuhOZUUGM70LPM/FK4zkkRmFLq9DtmZxPMkoc+cGjZDQOCXsA5tuV2Oh
NARax7VmOfXt7+46lkuZSTYx6b6EJr/l2cVzbq3VQSDDzDWqXnFlspONvEO308Mt
kpZYH9cEUoIOuVAK4HNwXkKDkWK9ynXA++dguv3UjmQwmbZqRpWUhKL/i2lo71dB
shQ4kQ/sNdBXJblhWJpYp/aW1+blO37vjTKWnfCFsT+IiuR9nJx7wjA0bnywZBF6
WZjd4pqCmEgFoYnpyHNgxGWek2at4j2ED5+r/hAaTZsULZFF4OtEzM7JAYGBLQH1
P6uF51yryJdYwFnqI3DgaTwT5jKYSIhkzoH0G8JjNZyKZUkChrjcMR22IOHVGoDC
vGD+t3mnu3iWZ1RUxYh7xvDz7a/nz51ndWLap+YHytZYqw23JTJv6bxmTKHYn8f0
Mhrs7W3fQx9TBRH/n3c+N1zGY+cH4FLgrKKF+LvzR1O4MhmvpdG1Lvhia4x5HLyp
duYI9dvBwAV+qoqnPMKTNK16zYqYDzf3LKj82jqz8SqjElUFCmyBvCvlMi9kWxDO
st/ZoBmyQeWanf4iElKh4Iss6TUKaOEtbs2EcDdk3uIvWsfmxF/JJjHClS3Q3ZkX
40SsxiIQG7DzJvYiORP8J7azDGnYo6jOff+j5Lc822c1nbHXOpTaByA2p5tG38kO
yTS7FGmL7ls9THGLmcyYHPKkNF6Nglamgilv3oCqg2fWyqMyxj5nj030ty7TCSvG
Aue9o+xcuxSuUu9ewd+Q06MgtdrPJbL3QsYmkiX6SpAADpr0/hVnlO6hOuOTD7tY
YlNJF6SGyDEQ6BAk49htSrswbccYCklep/2ywWC+mg58lCadlEFZ+wnAeS5x/LIo
8NMIvJrtho4mNqe3UgNjvEVjR6hCuE6EPs/fKwF7tpRdBdHb+4qxEA3Hry6M80Dr
zCWvSjcd38vsF+ilKSGZp6w/hoQaw6P1necoCdVvat9mHLcVdoOj2yHaA2eEeE6Y
p7BoLfxPrFraxIkLZb7x5rwPEWJ5oUuRaI4/Evm27FA6In++M95SiV3sI15NRd3f
vGyB5G2EBSJJgp14B9K3CXx1GKoT/++LyEFNVfVjtW1jHnwDsDQpj0UKb7IdSAYn
sYPSY0ub8GTcvOqJFpF+tYL6jQPkKAREmTSDSyuQVmhNhtd6XPJTat2PdOeKmOay
+zjhtJTajRyq3sxqYM8nTc7TxXvWvcu5jNbapXzoS0PhyQMNjpDYuLcu3KyQVnRI
g/VsIxWnIuC2KJg1SBAsTfdcIzTRUWoGgeZkdcKR7tP2KE9H9MejH3zVYuCzdNMI
nEdDGwPnV+Py2SViDKYhls1f8QoEomOXIPqppMiXRpVeb3a6tAoPbTc8Fz+rzM+W
MUCZpPFNlhiulvhJFbuhV/TUJA9nw0kY0mAhAXxrHE+sHl7Spei1EjdNue6sACNv
OYZhwS6Ig4CC+Tkj/BlyH2XV2f91c9HqXm5oPRfz5+SEWrcdxSiD4DCC3LKosUM3
EpQHaU3pIM334EsrPNZYpyqYXzoG6V4/wicuLysqrCgW1wEr1Ywj0lYGcWI3xdjJ
haLhTwpGbqy8A6rSScRqpcb7YvsWwk2SID0Gr3J7Vw+LCy2mDDHEgSVwnrA7Ac2J
KAryo7aofOgDwvbgC6yNQnXrqyyv0UZlGP3pEhQ5aQvKDz9BCt2IlKsJqnUUoq5h
H94rSHqdYx0eYU3iM/2Sd+faW1hny3pTxuZBcwWc3ZKDrC7fUMy2u7sns4B1xg7C
kRJfv1Rx2NhOKg5TwDWsGaXhZGSNLlVQ3RIoMD1/1ImXEPPWTSt38HYXuK6264cH
SgrePHzO4xMdafojfX9YlBfwzR1i8LRMFgxVflTBbuPQ3Ag/eFOtWZJwgRkUrsc1
99aAXYKf/n+9JYrdI0KYyRgjeVLDANiPpF42v3FK+dsA/Br+qFikWUN1rHCO9+qV
6PQterH9PxTf2lhE/5c8lOdJ6ogrWA6SgYlDxYpj3Lh35uA7Usp9cYQ5Z+qibYlH
7k3Kw430awYneOagW2O/mmHAgfK4Oi96dM1V/Ay+2RbZxG4dYpI3SN44ceHJrGVV
Xx7gL2VT50L/FZpl3TRKQqZov2rjHRps0DPmZM2vOLgGtxft7ygNFIDjuA/F3vUH
D4eevKuaOsMwLW76RgB/UlPMMiSh1O2eBEQsRhb7I/ctYftIcPrAKu+S4NJSaomQ
A7dkFi8X0ZwpGUq/9PAqREpDUR4CUJ/qDE3GIT2vx1LpmcEudLpUbG8LSDXRBBW9
6oxDhBTIumm2NOyelHsZjNog8opUuE/mmb+Xg0hYjVdJM2fuNRwctcs7pUR/TMH0
fsaapgnCGpWHNo/kXjr90fQTtZh/U96LWYmWWMWQ3oTdiWr4iTmtRZGMGhs/mu64
ktwWWyuc5fN4zFtMV3kp9a6yKCzInNPyoAuO2taqE1Zl5T/gMDaXnkxDv1qe0TZj
8NSJWyKZzidh6EQOZ9iSUMgEwJB0zuYtbIG/KMtmPLhPGj9d1DHCw/VE+JMrtUXH
xQS46V5BUEQ0dQR0mcAApHgliiSdYVjg3XIFNZ956wUbttAMK7bowdQ1L4sHCh3W
LUn2NgKage2Iw02CAlIsWU3tJkgJ5zFzuMw31NgnqUkGFEdzEzCWhLa5LCWtGx7w
yzW+Q8cBPXYwQcut27B0VxYvz1KschrqkZ/LW7utOp5zxGINgAcNf00D8IpGKujG
GnR6rl9bxCsCyD8DpVih8NUEXC5z+Dt4xz6dHohPvIF0poeHXXpUv6RmRT26Up8B
w520hE3MzAPUs/5ZhP7QAJF/i1LqkMe2025tln2chGMdj3q2QIwmPE+tIDKgtJdL
IeOo8XOlEjrLeXMMMNz62GiWTtDdq1kyVO57E9HF88Q4zNz/7yQOrmXDqf0rY8+4
kv74AJFXHxugfebWyW3fm0h0PJKhMG3RULOrQYLRUYpKYKyud/yRMfDjnx7H4pXW
XfcjEZjNRHP4l+Mw080Jhee6DNU3CkkDoSYg4Ig0m7tPJ6xVAk3o+QnGSEMxep9e
uXJcjvIpX9I7+C1it/j5BxJM9mKQKlShpifLPJDIPoLEqoMx6g/aUDlzMMDowLg4
SdM7+H/QB/O7TJr0kWsKFHgZHU0jrd5l0q5uVF7MsMR5/VpgOSxBJpes6ACEh79O
Q9UkZy8gQgmfYI0jaQd8DLeLjmmvwliH0hIER9U6FPUeJZx0gAq2OTIrmRseyq+X
Q5GZUT3Kt52UEyn454eFRb0vv6WCWy8+VxHiupwNIuvt3Tvq2pOeHPtXynIJdoey
zD4XVaV5RSzH34Dgdsnnn/xFHC7nJer0v7GaPP7RsDd+nqa6U0vND3j1FQ/UICoq
UUosrdxDLEGB867cu6fb1Qnf6V57lHuLIo+71nZyKpYdrxUmw/iQzMQalw3kZ/Oz
zToYRY3Oz4H8D1XEWtqh9ZxQml93OKbOPJOTE/2/DvLOZLMBhlo60rCsGj0GxrBy
ebJ3AH2ufuHJqB6yUjHiO2wLlBhPZXwcqOwp7q19JnIlXuq78uthlLpBSSNPpKDg
50GYFXBrclpGAEbxXVXpplSw0SZXI3oyhOMUMtgd5o8jHwXI1AbHuF7/1AZozwQP
bRMO+uvtAFztFemuIbL+1c+CWRtoo9rlBMbpK7GAs/ezRgv0bYHcT9Hdtatrr8Ic
Ggs0+i87sTz9rxYyU/NtLT3OaoEEEXSEBLrdxCzbjPvPlPRBcAYiQOHLum3b7gmE
asgX6NeewfWdULgT9D1cZhhqJgaF39GJx2vLGqGtMZKjXe2Mfxx8b69fEYlL5fMB
7vMrA2QkCJPoc4wN564dsQneQ7UnZH/JNB/UCpDKOtoB2l+xLlBh9LOwGlIynx/N
tgGsd7UaHHaYBTQg7auLnyLKd2fYgGd5qKyEvJfmC/jy3JaxlhzxefnQMi4QbzJu
EN5Y8NgewiIow/HbDo1U3aKYNq7v8xShN5hjqAreWDcus2N8T5lhZi4jH3ys69Vh
swXq1TyX7FoIvbU9eWJ1ZEcutR4wekI2ad+26KNSBdEQmhFIo6/0/NllDodVjg7P
Qq3uObs7yrkaGiEcgfq0zfamwvCJuSKr31cQMIEzNl+O0yGLQzXGbA92FL7rzeWF
4rOb/lcBPNXZrXx7g1xJRPZ+yLNuWD587OsIlYKsViAK+eIc9qe+129eFyGyTufx
Ew0pJGPom6s3+Gr6o0fvqrD9yT3sjSbyVV8e4WWoB9yoEK7Gpa6TbwrsBwQ5dGAV
fZ8NgIROuMGg5UNvzbf5FM/DUo1xzMApNRo1BuJxv/BwUKie9nq9HCGHGjxHsVH1
oacqRbZ/ICiZBLpnRJg2g3A0XO8sa66y3mFf0Dm05O5HRSdCO1Db5v8p811/WRG2
+IpkhFZTOlRa0SnEyb/z/vjXijLAcZt37RfRisnJ/0kH42iGm/57fSGB14fxDNwQ
xg5bEZmxeBpPIRUwr0fB5EsLXZZMQHYteIKndpMlt7phnVs9sdpDLnmBNLbxg1JV
KS39K05FfkFnDBF3oVVahnawsnqDXN+MrnVroxKNHmx4V0W6wkJWHREJBqSUmr+0
LSyP7ney8bPdAao+KmHn7I7XQ++o1ScWhp25PmaqjkdnnTUnBkOmQLi81RzTNuFy
I7thLVDO27AYBy2BGJ6+mNYw/ZBNvYjMfulu189wbyMscy732GXQpTGMBBn0rlCg
HbbDiYHU/SNwaM6CfpFf3wh+d4DtiptvdXmu6LzR2Q61EPuhrTzHzU19l1Mw13xE
67ACHEGwCuHfXkEvzo1L/TQhk3cmGzw4WH77hYF4f4obsnVPJeYIU/HpqZ9HOPFt
GHSI6Vgr9zt2kFHTlEx+D+HlR+6kv3pRyeK/050VbOjlU4wMp1RUhwWJ0iQWx72Y
hfxoacNqfseiyL40dfZ/W0tmuOmGJPHOQfSCcnfJcfLOpwR+U4RNvK6a/UpwaIuu
X1bpvU5FgiqRG7t+eo50lbF2xTUSfgtdFrvaWSmymR4EcNOTxMyRj6VesQDAes8n
zgHrbPnY3G4KgzNWoQBXyfU5s7WqP86hHzh8jZ0SD5cpBSpsq87Na/ARC1Lc8eKa
Hxb021rbk7pIigTmOQD6b95nIXMWGC6hSncno+E5wlA0Ol0Fu56gQ3s3/vQ77rM0
sG8xMI5LukJJPRqzK4QPVV5dAzG6aCtRu9QpYHusUgRqBCqvFkXCgS/QAZ2eB04k
PrVKidDiCPa8MVuayz453PCNx1jM+ZexjBS1kYVN5SKF7NtjgIK+ODV7YRJqvjcb
XMBH0ce7va5Hrk44AABADPlLVaGh5z/4TYso3Jv7uiK7w0JQi6RiXRahc9UQ9U0x
eKfr2/S+G8JTcmOukxtU+m1Jqv8dRHUgwae7nY+1K+YpnNIKJYeGSe3orTpC6ROS
VzkD56L/37Wg6napkbcIcOgTUiutpvUN/NSoe3oMfgRPvVlOGwUF35aWhk6Ovyf2
yfsDZ8iPXWxT0coHUx1Osg1QAfdEx9jslZf87PcojQI/8hNdFWgAj+oRv4TK3nKA
wN6ATIMfPEk7Nmcj4SGgDtrWOzw8strijLq0B6u7wdz5lQCqyP3xdQ/qWRATfg4+
nti4MKSUXshbC2o5+cyCDKmYgtu6KIfRZE357rjz/YeqrNvbY0w9+9Gt+ON8Kqpz
Oc5AIIeRw6oPdnbor00kg7Tl853HaIuizp1I/bd2magcojFAgOyunQBO7So28JxB
UJ3QB3WiiFeDarhDUk0cDxoqa+D3Ojw+SCxQPqLiK5vut5nvn347SnTdkqhkBjfl
GTQRq6rlp89RBu5VQT5NEM2XZAyqhnpMutYeqABdUIspfCe4fXmEeUddkdbLAAf2
K6Ea1PFznC5uNqGEN2eM7GCQHqkt6kZvBHt4TOSms+UfFj6WnxzW4eW2D3OSDLh6
h5eRNzBiBBuqB5RKsBT4nr64aDqg85atKx7m5vVNjJ1sCJr9mVQRNFh6gbzxFlcQ
qRhY2S9YfPpCfXf7VKhIHyg4luP56HozEAi64WaFxwExcsZeqEI6u2HYHUJ8pCX6
Odza//DlQDgoPN3AOlWextyPZQ58TBVHbvVxY31O+O6LFj51y2Ek7fVhIIYjINRi
jEPe7X+Qiyj44/0JKSIjmchEUqeeWvv/AdGScirKkzJL/SIdNaqvp/0CtFaQY0T+
r+fHlFgZbR0AJ6WcSbWI36cHqQcBHZ6pSH5Uybie7y7ZcvNjwJyG2AMHw/4cRVYK
w+FIaxuS153wXxxNKGYkMmLl1GVBeSVBkq2Khp7LHoiBRTV8FgRlbYQBMsm3QP2A
d1mjTME27ft+ulTS2gXTZVijowc5aHsUym9HC6r8eFMEPHUMOjjQ5/396cdiv1D5
GtWG3pGcjBDswqDc+G47xe08iMzM8HDXiqoxUVZn7P3slIs8l/QxMBr5p516zxPQ
bsgRVKz54qQl14q0m+puDTYN00stqQUb1LKOVotT7os4BdgzvIYXldrFRVgcOP/8
0ivbYG2C+i9TBmvTW2VWKuQSUjU6Yz8/WRmTf7gQJ6cpO7BgdvYgRumvM5gCOX6g
pY0qhXbNQj6+lLk47K4Zf0UQL4JO2ZWoiPEdI3y9GiRJlD0g1enTHM80g/g6YLtI
rp7np8xngATwae7TXQAbZWkZhumWTcLv9wsW0xZbDHZegjYQ/3LzVhW1Q0EYyiV4
LLuCGX6xCrnqZD1L1l7JJdDaCKCwkglBY8zj0Y/h2eSjkkJx4/yRic+QF0zHcWpb
PpoO3uUcSY3selm7UDfbzakb90RaptUV7u3LshSEgCFJKRD2+Vc8NWBaQLuDmdTL
sJyhH8xqLCFgjQ79h2rJ6Em7NHqzeoiBsUjaeD2bwUrW8pbLhcB3rt+WbKbXZtlS
D+192eM/yJioG0Pe0LwcBdphaqqeynmNTVcLaOAsB/Mrf9hC1RegOkGKqlp1l1tS
hAGeluCNLIx/7u1JnWirapJFNsgfepTplF3RMEUPPQ71aqYTN+LLxzO227YzuyPC
fHUj/Eb123sjA26HVysqgqwPrEVxvjpmYNya8c3iUYw9Whcd6puXzG2N9OC1LSyv
n6pwVo7lKAbyzYsk6TNIKc/Cynv6P+tyH6UrLFKI/Yldvfo5BF+zlKInkBzCfKEi
0TSm4ZA7oYIbLAwDqWZ6uvJuqEYqIbyEHO6NnTOrbDGU6MBvTzYpZx/vDvrFOq+b
9CWr+1aB/Yv3c/8P3YY4SmG6l+g7zfZ+Tg+Y/xq/NnjH8EpjS9eB0gNfVO9z4cUE
shg1utTcxV/hGIbcVRov/NX7Hsq3WIXsj7YEjmfWMrJ4Yph6kp9jUT6an7UP3te7
bWy57I5lQ1bu6bo8MUuVgg+cA/G5Ko9SUG/iHUx9KaP7SCAv/A/RnHmXovnfU2Ck
Hemou2N+Pf0tfmtdpxrvf9j0mV8+2dFxu3Js5ar6ki1Z17m0yW1F1RHlGMnTXRZm
B6uMu+JOUjCgIL+27hLUgRzbQ6rIsn3pgMfn0nfeO7VBCwZYh3YvHbXysVlB+NaT
fgAGsZQQHTAGAWFXNuGzocRoIwvgWmTYVzNrrS6y71yP2iVWbjBu3rkXtb18mz9V
axKTz93XRiefPQgZmyCH2uUQNX/HnTlXqHkl8j29S/+q8FOaV/nvxPuinAE44kzh
YwDQPZ0PhDvSzwyvVpstpVXaYd9V1AFZZQjS7OzsTGWhr/Udi4eooGDGuY2XJH8n
DbJSJU3FyMDIqzhoFPIjr2Ic68wALbqaRchbaJ0VguHdLmh6WW2y1OFRZCpzvxaH
Vwz0qXwPfgBd/sDWzhpPlDQuikXN63tM7m0VFE9xUQmwGMRUTmLghz7uroo2C8nE
crvFBRGIXulQnKOLuc98m5lD9qwUdhR6O/+eIRFe8Myq6J+LNvqbDCf4i04XhTT4
Uj96xbxs6ScAC3DCGOhk5i8kwfmqHtVXRldeMKIzYfik4TsHIHinAjCFlAUEfs+R
26Aar+j4gFZYoG/2TfIii1Kd55ArMu4nzCgww/XqoMWutGG11omdbc9lgen08UDO
VdLILej32g/Nw8bsNOBGLapZ/t/Sp4BNyrTVVQWTsAkioXJRmjvkWpUYq6aHjfdX
fqJnE3xrPlkdw9bx61xYxTn0PgTZRS1wYA9kPBJ0zqUTE3WRPHGGXpbh/XokEiLk
ZPuQUzA//UpwS3ABbhvUBp+OJldrkz+g4M/PV0vtCWbGVva2/DCCLeKorIAalkP5
mDsQblsVCq3SV8CClD32OYCWX7EwfKsAiyQgg1ZxZYCa+74j4Io3oqJNqQw9qtg/
1MM074Yw0P74aKAQnmlidGwN4+8CD1HTJbLb5rL2P5GVPIRHDVAPDUCe1/auEG2k
Zibf88PI6hePKv86pGYVqRCvmVTwnsXwUZ6Wm96lMdCY27UoZFSrv3nPwxGnSiSX
4i6ACNY3fWO/PtTjU8m3SPKCRc3IXnhN3JkePEyPdujRecOY/4kCq8djp84IxyEK
qDjAux8wAuF5kRYV506sQf2OR95/VHqZWwzUrsXUD41zkIm1ghuyV1O7G95QQSSE
4ljRNVSU8HxCeJW8CPILFw8fBlDqVbhuC+J8r8/VuWtGpqD9D1FtL1UcE3TlEqI2
wQDDa45C3r0XzGS+Llx4BrTaQxDsKPyMBjgxgUOsrp0mV1AcU/A2ai+MMZuzklvT
5V6WXtk0w1kKMHBlQ8ubSRLIJul1JYbhAVLID8/Pe+JOnuscz6NpkAOLu9qaGv4K
YyJPScpTyZsIn3dPdOvFw0bqQy0rvsCMK4D4959TeJCtoYLvN6UQDM4r51nqeAxD
iBR5OYHGLbNw83tuErLwGXCwXFtH3mZ3G0fzNMMc5bhBW5t6zJ3+HUyBRyZxE5l1
+SrdISPiADEFX0CD31ydCEsjtidH4uvhK3zALuxGQ0ARU3/1OvSna1ZdnEy2xF6O
ZJBcvNDeA1bkaSzO6yLhKwzask5xZCU1JT2RPxdzA1pRD2NUde4d/Hc17n/Cr96S
5GLeOE8AMMeMUgkleuxd/b4tFYH7+M9cH6GbPUHHbvRuAxoKrhkKvB1Hfp2DmQjL
RDV5YESbPQAoMRxUc9biPFAyUbpi5k1IDUvp61upcE12Z7zmm9CHtqIpXS1SA99U
M7mSlK37xVYoXQPNQkjdnkjsofd5yD+IpveP3xguL4HJ3/hl96BosD4oTldupICs
9GL97GBtpZNyF3M1lsclEkdM/xPDnyCP5efsTsQjq3Ivpg6ugTsBtf++veUmwS9Y
/bXseqhiispTNHl3q4c4iKqwHgLIqnY1KzHZzIAzoOcGWI6ZPFNzoUhHnpUXk1Y9
76yJn1T0se2E2+PxA6ujQ/MSyuSYd7Y/8y38ROxjEnqKr3kHCQMoz3k8dOJTM3f5
RGqhEWY3KEHTKqydTw+9ny1f2VFCuXL61e1wlvKZo23WelmTsBRgoWm7kk++4a7b
d7VYiEDypY323fxsZ9PvA5nfxjKHh9TpjO1eVBo/QvJBrUOvb8Xq/707FmnDHuUt
XBW4ADE7/1X5m+pPL7bsIXo6raGEaNi9oC156DoK95LA2TOgOoEbVYLzof1C2H9K
z3/MVdcosqsNT5i3ePa1raoUWbsqlu/bPkY0z0+eU0kx8nk0f+lzBrNeVow7M5Tl
EPM0PDQW7CZvhgO0qjl0h55b6rTQMdOFb+X978E0HIXoXpEjhtrVzjU36R8EH/8+
wFFHMmLEvuiBrtiV34QRd2eMQtvttyJ19dWLMF/mLEXGvvaeltM4cNR0q88Z0/VV
mGCN661mqdROzKknHdDLxEU6LAyQnadlFWi+ByEd9Im5IcLu5hkQtM6DtvyqtBez
AudwnDTsh6Yllul1zy1qvhoRQe43f1RH0mzDp2W2C9gJo+Ynxhcf2KUuwFePkmEC
8MEqXUFqdM3H9KHHeE/GZeMLc7JXfVSz23SLARHZeuzwO1iTbLsZ5tkWLv6I5vcG
U3veFeU/sbzyDv3if/zhURwIRC/5foHOuZi80pNTNvIjRQ9jnYcSyXtLezrX5c44
Lv2B7G/adOF+j13ZypQQscNdc4K3nwLIm3BI5E84dTPf0WO1CLqZPP+MDnvH4xCG
iqFy0CkSf/fvqVWK+g19eF+MdCJlhdJmsBptO+rVpt4zP4InsCtRJ6YKGmxmdrRP
Ojnm17SRBQVpUT5HHkJ1SPerJYESd+pXBrvCxdd2mgBIpKiaP6i/HqhK3I7FIhU+
0/vI5ggH0exffAO1S4yW/b/jgNN457v3LN0x3DxLD9jFQTWgLVXzDYLKTg7HQBHB
z3aT6yNVY2QNVrruYYDNDLKrYvwEClj+HPC5MlH5t3RnohHyM/eANTAQVN1r+IwS
V6oWlWdLSBaw7bEDXRCfQt8FUsH37k1xJsTgrjpdQlBCFJ5nSo/fhxynP929UESK
s+3sRnp6+rVC8VBnxbmLmpbDoe6VUTqzEnngdZkhfT9zXot5Q37wfk/qGRM7Xaw3
YvetKEJm8TPicNfRjNlXeo09qxVZygcVjb23NJgWKwsmN/7V4P0+V86lrTtIEoM1
MqiRhNHatIRRcsoYTLhszDCm2l+vA2y6X6tZSYsGu4VoY8Zjd7GPKHIrgXAiZ0+y
2mj+t+QPZh8d8kT+1c26SdpxVRZf8Ax8KOMhL2d7wLgyXxB3hqbjNn5ttTgP0iIh
ZBK4yxQ+aqxb61lvSC9qrfjAOnBrEzfFkHFmEToqLsvBTD0Z2exvw3Mb8qyk7EGz
UTBocirOuFyFDd1ilzfNQFpWYZb0izb8R1ZjVceOMJFus99qJWQVQigL2xLwIA+m
SiV7FsGaXTxiuInbGlBxY0ufGUcyJlxXtBkrxSPRTpcURY+XU5njNCh8NMJzWulO
R8EDsiKpRnHnaRCm6zqV5c0LZz4YP5GcKV4EEcAuaqicCauDuxyPu0bf5ChJ1D58
2QgNKOy4KouqC3HIRtfAxoPvlzfIz706wf3FhdYEPGtVvAQW4VnCW7XBb/LbW/l4
RzdziAhD0Ubq4RRVeUNcKQMMN7OQFRdR4C43iXEIcjes7OMwCz6QVzEe+bsJh2LW
7/40f7rjrw/c/mEIVFaxOsVFmSQipXJolk3eRSfuXQgv6PAeLoNYTJU/2oDP+4yt
vVwo/KUM/bgKKMM6mpvOwY5AyB45hsu/ZpL1DEv3Tm4b10+dggH+152KI2D1iqfn
2rzef/LlD4bDgTwmfMtQPmnI2G8XBPQT394iLgyElQLznykxE6SyIM0JEXE/husG
8VNrpsZ60t6p7Dc3GXOJjB7ehOaP9RkpGxw3s5P99v31zZn7l5xUtY7Dmvgy/gjf
pYT2pKDD9/oviftwtGGutrqzcrOozJzkcwFuToMqkljIEpvhWeBfgjedVuitrKEe
ayUcdUn3JNI7UkedtzNkbOmZDll15He5rajoffMBLBFMwgpEWsISZ028SkbyLL4A
sISnxFaQg2+68qfKgJGfBxaWWMrL/sCr/jORKfC/ePURrIYGm5bEmfGS+Kq4FHQ6
JIZFv4FGjcg7xKB8onLluQytKW0srXFWO7CKaWdY2pUilA05eeKq0MpjsoS8Q6k4
9hecxYIDrKjm+P/v4ysg7ylESuSUfYXmkU6wt74LsCANVddKwB3HSraqkhr6K/lM
M8Nop16JODKZcn3+iqu2jC0XdG596Qn0WLW5N26OhGq1caWfhfdBT88O+lfZfHE6
LTznbiZi63Rq2EEIvNAb7LapSUSgyb9FF6xNNu5jgEqWmmrGjA807WLmKqdhMNUv
jrcV9/AedfiwvT/8xymjzPnjxxXowX8cLLcK9PN+FYWwMYHPqdlY3F3e/4G9xuG/
km3o8fltafXt7UVGgaz0r2Y1UA5ub3vH8sewv8TjRSvkyZCbpCh/FTqgFAArHzwC
pULlgStFdbc0+6gkz4j48n/ZH0Kmcy6wZ5vG8FGfAViI71xD+HKwjz5Rfx2fM3A6
7W9BskpsHtDkbReeA9hVgeBX9dFsLu8fsbTo/+ZYpRsGDi3XZypoicGG7lpnzMQj
5jyimw3kBvcyVUE3Vg41KpnxAAl6tTDhQv5TM00TqraqDkO1wd12C8XXPDoHSKLW
5BpeN7YkRYtebYIHjMl+WUZQcLEk02Co+qJ/W5YOpwcv5FpNSz3xJqkKQyZ1Tmi7
55igMDhJej2xRhnkA0UMwv1MCaI4+nCrmGFmXcNszE2WNbqedJJhhVbAOsN+W7pN
ZFiOlTlJ55EbaVAvwZbZfUsN0CZk5NhfmgTvlA25lSdhCYYij5xHKEbB4/h7XgN5
mrgDkJ8p4il+psRCFrHkQAQKaPnq766j76nfY6QR33zV1soDT0e0ETW0XMp8rA5Z
l5lEe5fdcXKERyCQ6zWAyBPR9XmE0w9NZlbwFVpaGSrVlFTAGW98rOa2IHZMjOxc
c5OGLTApsFthdOd0VM6AuEAxKunuTc1UwGjVOBNKRGTD/wzjAIwUYMKEwm5CaIq2
voZxItHZi6rajDwH8WB40pl3HjBrXJkm/pxXRA4JS18xnCn0KFcp5XmQGHAXJql7
g7+qie/EPlruyqh+mjXuCwPDEZvueP9P0na0isI78NvovQMAZjOL+QJBqurisjBj
G3qN1cL/3uaPUoYqL/9xkqD9mY/pgBKG1vbLnoQqGNiuFrvfmn5OSy4M4RY8ZxZF
AxnDacEsY6wF0IqsJnBEi0YO4GN22CcHA2wSb1FGSNHW3PJvwGgyP4ya50aP0o/q
7jMrqTZQqrG5E0dbUeYWfV9nkj79xNJNFvLcYz2wQCDlfx7NvJiPFvPxqmTpC+r/
iaUIwIVi2vKNaR8kiCPvuKOn0x5/10H4axjO1t3zELjLQ21pzG4ydJ+Rxck2kWD0
+gt84mMNTXQhpIMA/lMy49hKtcqLqRqaIehtU1bcnwwUAqghj5seUmiDGa+lRmYZ
AbJVakwKsI3Wfv/hh6655xwOIsIL5XtBbyWnCdEOZFntYruf9I05Ut936zPwmktf
tSvCSvWb0csvMdKNsiTDRcQZAKu2PDCwkgDPDNilonuoE13VNI9Xa8NQD9xVxluu
FOHwa+gFIfMLdpcdIB1eGPDpZUn+fvKn5TqdBD+cG+k2/ZEc0M0U137Mfm+BJD9t
2XAjiVVKVPXtCHSDibuWHGRFEUmOJgA6T9FUtGeeF/asugb8MVNkTIC5Q4qnEv9i
WTmywd6AlayyEFNPtRssBAOQ3hEmyXx8hHLUABSkd+IoBYuVAoa5oUda8B97MuiT
bhg8oKPWbvEnP9Q85nk1x0GB6a84voUCLPHU4LxfY6TPNV9fNQ9e8uQYolh/hpLF
gp7a5058AZMyotfjI9MzY6eXUQsDlBAVV3URL/tU9IvaDjRKKZaQANYGfY7Iifb6
WpbuZ67SxZe6jHC+M5XO4oR9hF1E4OEkM8INQQRx5xs28o77khi1LP+0at92gcO5
GZ5ReiS+1PoEpC3mjCPp29JUePb53IvsGIqfYU1cLaRvfTM5n8FExv1efY0imRQ3
q1zz0idZNl8AvSM5NRgfKfoMe+ziQ7IErjGlLK3QpqM19prXyZsOhJD3VU+cgaHF
9Smdp7q++OaOW5F4NMQS6e+iOIBi6nrWuo0AzjqVhOHRZPBcNkmH62jwu8FLk9FV
GNbp/60JzOJtpokZrQc8QgpxsmHqnsKeF4HriG1654pBkeQpkR5eaNonHrByhpj/
+JBpEx5OtZWXPKEEg3dF10fB06fj6zERMBZkoQQQrkwgU2MYbSOLuNUU0+XWrwC+
J02Pj1SawZHfiNhiErEGDRvAnCAHV/h5DsVaBnPqNzivyLaRMsn4+nZVq6RTh289
/VAJzxuHnVqBHJFuy1Fg8lxc646qMNepAR7XoFupYPEkw2GRN9bLBllfkUSCWpmW
KKapBn1hVAvKZK4QFwmdJdB2ZR4MWFlyUVucgrDZb2t3BP3eksFkC3grAVSrxeAX
qs9b9L4H6G0c/vsJw6y85aTNxLpagHVQvneQw3Oalqh9GcwVuAHQ9Of9qIqEFzqF
bXUF2z0NFs9fwscduGBbHAJ8OUch15mHJ+0xleQqC996EZkI959FhSGdQ8QQRh2c
vn34E7F2OW0XzASSWgu7oqkH+b5sp1LplhkB/JXfMk2o2g9Qp3wR5nmfxtaDkvMs
rZlAt1icP0qLWGpDBnVt9M6+PjKy9hk9kYiFi0jnqOxV9CUpd1bLiZUnzWgDkGUJ
aNg+AkJjhjbQV1e2Sqe63/K/gTZI/9flY4wQ7XK/ytF+dwxtMYn/R2EP5MjcFKMa
nbDFsL95dA8lMtnP+AOruJCh4HLe/f0lYOW3aggb8XgPRMYL1nxMPJRJsrPM4gDZ
UBotEKc+t6nNDpc3F0bqozDOkcEgRDBDA+U2zmzuMQC3ux+5vdNMvXhvRlBYv0I5
Yvie+Q03XFcYOoSqv5TVzWfC6ZiMdNykdUZ0VXAd9AGRBHB2Yb7kmMktflXHItUA
zq1/+zfcMMHZYgyNm9TYKEyWdn1GaPDFsob8yerS0d9ltE3RHNCfknanIE3q+D6+
BZM4IW6AOG5NDsSIGGvFVUWZYVKVRyRl431/V9GComMyRP4nclwT32mUsaDKZKfx
A0GOAsw29xWy22dTuEBuRAT2em3pXUBV3YggOkDXvJRK+z2voAOTEnFmjeLvS8qT
cSPdkLbFKdRiRi3VTC65EqsnNh1TA8w3BEfiL9nrmyOEGIeJzeZicH0sQ8rw46j3
i29jF3BIoyG4yf6j/Tjkgh/FGayITsi92emxUMufqiW56gmeXGVnd6oPW1OoBxIi
A+n6/PX/+WF6iFMN0AViByiZtngdi5ekUnrOKxJ9cM3Ti1a4s/ZcZWEhK3Hk/6Ph
qTJi3e5xtsYvrmCDjiQpAwKHbj2rSoVYDc99K4IQaWEabJXod8F9/hIG7YPJAKx6
HYCtk5PhnMDEGwhbG+yWr9ic3O48j+UiCcenmVjSnT1UPhmhLno0OrlxjjyjJymp
oR7N8kzNqZSR8X+ycMW7+ybMh/jKd111P42cVxR+170+RsxTILlxhXQO4aMntAic
NexRvyOR/4B8TKZoeJvFF09lQMr/+FricPWYHzshZcDr7dyab2hrFhgfJEGwX1yD
LkIAJg4+ZIvDIeh6xG8QB/omSltdcTtHx/wIgr3WP8Fs6L0F59DUlqfLm2uoovXS
J2L/ShjgnLruh28035h98YMJan1rdh5TUoVhJSzPJXRxU28fOK0eKXFSd2dGYWoL
HVbL2/3wCAZ+NxgI3vdXdB1LwzwUm302qgyUeyLzZu+AaMin4gSVj9UvxZ9A0DHm
f6FNC85Py0fOg8doObbCgKIPs1J0aFZSNWATe2XC1S4ew3fiBqVGiq3sUJBzy5Fl
+ES5INt1X2HYUVzYjf6oelmRMcb7kGCBJauMcpYeVpsSVDPntlrcm/i4NjRK2XJR
iPbvX6gPIKggzOct/eyFMHT1qgOaa63iJ/cxVvNoWI+BFpM2YVZPAdRilgxzw3Ex
YjFILr7cZ4wMgaUKeFNFvkRleeV1OE1sZTrT++3XMDaNj6amKowiqHxwdGcCP6Tp
EDD7YAaBpDSHfAPHqdX1FbZjPY+qbcDufFEcvR3ZUsoSsQh5n4GZXk8m4E1G43jD
xKXIA0NnZPqYat/nNs+H62QNQNVEUDT8qn7QW/HHeBf0hllycVmvkZChAEp+LVeS
1o8KO4fgfRR3vgXdJI/JrCKT9wfaeMnAkurGBhu92v2p3lKwlOYPSLvNk/2ZUQPc
L9UGSHjwD4lNqStTi8zCrnxlXBcPWdzgAb0eOyN1I2DesWfPi8PR2xz4Uil9UlKU
5OCYUsHUgW5T+Lk8/G0iwwBqZKnjtQs8aFwoMDBDLGffqbh3FlrCYjUXBtNzC6AP
L5A1cjPHQQTq0fQp0pm6FiSg3hPFgP28eNxu1HNqc5n2zZzYC9tzEtcxGBoGaoGo
pIeTMqtEqCuGbmypSKvybOe7MebyDtXxlo6jl7dnMN5xNkuMh4IZalDSmD0mZu5M
A14ndABI+ZNmTHjF1b/gHienEHTHfYv9NCUcpIm8BaiVC4cmITwQgpdnjgg90ouz
yF1cfHqqmxKRNulalBlS6xub2rJkgAwt/lxaXbmnBFO2obs/POxa710DJevwLbUc
1ePFLEfSITMD6IKE1gZQYsWX4q+fTp7s3R75Q9RvGTXNxb2MmP6HUleto8bWCEGt
HgLq/QOv3xBegfOLbiBZoStjA7OjgpC9e5WYJPyy6hppbN+PalYOuS/r8E+gAs3n
f4IiRXjhj57azM9Trl96zmuQzLgdCHJNb9nRDfY/zTzmP1gze6LGtBVq3+oW5kfp
R4MIGfFCSMfepvL1/Fn/l34941JIfIGhmCWhJ4QxwTVpFGUdLmDa9lzABRqvE+0R
MRvTOcgA99Vt/W/9jF2ww+j6XRb7f4NTUWmML4a836JVv8u/rsnWu7RdnrEnjEcA
bC8YMYs5qT1XbTHd/s779dEq+TK3AGeyuW52JimLiDNej3FhXcUc0CZqRViql0YC
KZjQwu3U4PhHN7bbaXj8bXQiIHY0eMR2zkrXhEzhKWvpl92uBiSBU2Lc9MCUfT6p
g90Q56yprYfEV4KQH7A6JH1K3MqkhWrrIULv47ZGKO9R1NbE39iNeKwuES0JqhY7
ottdCxSF2KxvCoYxuPzq6trTLTynw8Anz/JmKrgqg7FkFirFWIsWS1LCn1KG12aX
i5ytmIoeuzeqcxCUFMcW8Q7kmOVS2MZgPL6bRpcQgbuwrPSpk1hi8mixKt+oEejZ
ogmnijrFfHRoYPriGwPk6u5bU9AwF5fkOtbSamSx3VZpbzC9JdZbKPyNJ4H8TYwR
TD+oxjjshdG2PnogvY3/ZMBecLNMznyg+fxTHhv+kW4mqwwj76lgdf+MNQEBkwJM
NLND4vikP3BjFWuawoakvl4Vs8QrzxKKgA6rp1osCyGQp073cCIHRN8EPCE6d6Kt
JOI497EQxsVBkRvP70lqml3xBgx68CpcoAYH+J7Vr2TofrmNILJg+ZqqnqYbaQKZ
+bKw4PA5aATISGfIWCNAvTdli+fImx+mEbhckNObwbWflP7w1XgyWebKdFxf84XE
PZseTQKwPLESAZKjzQ0qIKilfcI4RB+ie6ngYSqdkYP5iXMp2Wu+MpxPPHzHGFIQ
GDlMIvsbS9uRP2gA2kQFCyQwSYU5WX6vatrZlf6h4N/YNrrr+VU5IJWj71iRmN18
VMjPd3hJCE4x1KQ1/97Dd40BK5rv0Y2EnEadK7pmkQWp+9/TE1uLOOrWrOMxyPTz
zbKJwQJHK8dbNQCkNzBGcCAvdbG91hHuKA8HMCb7SuKp556yVAoA7Ec8weh/MuVd
pRE7Hd7u5bzOGI9wFDaMYjxG44GgfDkJq01yg2w8yQXFz6xVUkTjkz28zcrVmvwz
jZPs86K5amhX5er1HKnfJVxx+cU2j95cA3vj1ykoC86ARal6KCtcO3bbhHDCX9sk
tJGVKRkrENAwTzhchjiONZGwF4uUb2A6/w5l7bQKRv1Pq1L+xVtxQbWYPDs5ak5V
c7OF9teM4KR55mZaYJzU79Qyh5u3S5s+R7KDBfwN/C+JSq8+sjQCs99usxIa+xWq
/JKqtnV822ThnbQx6UKDcmrlgWNe7PLAqZg4/O4c/mGNqhlxF8k2Ue+Hfgw9lgrL
b2XY4/exPDdiHYi6t99zQjiFt7CxMUGrl5RlpC5itO16fTx0z171ya+UNCbjzENv
1Me5TG/3VOOdLwC6He6V4y+B0BI0dRyj6y5n3grTaHMQZN3Kn0JCbd0vZQ00LduA
Caul9Q46PaVwv7yf7qzLz3Q+oY/GHJCP4yj30ZqK/kYMJTgdSLSzNXLAsyzaZg+c
MgEc73N82uY4nKBFi4+AnIPX2wPgRBf3MiiGF18G0YoAD0fon/cdqYH9mntfzn43
DDO/q2xC2ZHerI3M0D1/k8v+4J9uhEkHl4wbmNpkSdvDJQCmRwHUwS0YYa1km2TT
/qJALunwTnfGJzwlyQJnP9fdDSmvoabqW2Iu/i26+TcL2oUd2duNhmbMPMpYB96P
M8cItYXW7i6/Dr3pd4gsT9Nw3Dufz175JemhNSdIak5b0GFvLaaRZ+u+cVAhOL/V
oL8q3xe497Yr6WdVOSNtJ1fFc6F8gn5hq6EDM4iW8kfFSGljwDP3yeDt0k0YK9Dk
YeSR0MGeogZlIkQHfLk9dutNNNS0Hj5s7XPVlMTKQBcqzo8XW0TjO7p2GbgcUui4
cfI6xnxDDYMIS7751vdbSjo3dqnmGcliqbtMykUQnj1v4pgPSzluDL+166XM+WIt
fFzlTEt2DqG/KQtwxx4xEOoTdQ/d/hwqDWVm2W2PBQG7Uam6AgvncWLNe41Z0yuW
m7mEg+su3qo4GbG7jHcH3i/jfmZQSM39Gl2Gv3ccKWMlPQ/vuxBCavQyrvWoDRIR
a/mPmoRYZxBtgVvCffggOP1rOERdE2u//5c6vfiFTFo7039/7/cpsbYLOfN9IAZG
z5np7c5AXpPImyDKW0iIzG73MvPdfsHQUY/K/YtUYM/H9j07WmKFpehAVw0f1Zjy
qE1L4UDT6Q0eJ28flGmApjvMJP3hQrJoGgm0ElqEjm/gg/RKwlwbtrTdqscbNeYv
OziMQVHRDSgUqqBiOyF51kWYVtx4m8dO5FVbJZ/1ibbrwRu8M9RzVrvrczV+64pR
H4hSvE9dLMQj16UC3XNsmpn5oZSQTpW2pMC0NlcgcET3/y7xfmq88hFMBjxNE3KI
TgUClGB6V/rRH45hA8BpkpVqYnGdlF1haWy3bf6tnCF+QJiu8qNzoPLFcn4lNrEp
z3ZweiRpTOPOSdKAzxAZSG4V/JZhBb8xXy12tajNDO5vPxvnTkmK3FFUhf8dno0S
6/0akH4ZBwex1SQfpJDEsawvAcdeSGpUEdXBPSJnltUXdELmijb8w6mO6dKJeRtY
04+43oNViQtKAMcB/W4DKYt7KEqTsJb5Fc0IDg+KIZYcDmj+N97Gy9iKagqU3kSi
B/qU/zFB7NyZJTJT/EdrrqxSSp5xYSDVeuPqQy4ZyMaXmOGRG4V0yJ8SUUpMUuOG
TcLboDXXJCka+Psin2OljZ2Jx98P70ELAHAKOwkegxspy9G05ydQe/313ci5015K
bv3VCbHP1FWDaKDOsXZpFRDa4HCeIME3+RDvWkmosPXItIEp3Co3HdaXQYMWJ45E
2bCgZE0/28ctT35J8q3i6USx+qY2FRjsXaGZ5xJ+cQzXelju8lLkBGhjLY7mXiFs
FTuTQwsA4r2bY8qHwdvS2uMyu/fKrOmu3TClla70gc5mPKv63j1VdV7PxtUfJsmm
zYF4U2Rb6+ea6/sfIT8aycFqsyD2ZessJfjd4AWCFt7kOgwwWnZ2kavPPS2isq90
8SpdD//Gyv13+F2Dq/AmAcnONdYtQu17ZwSWSrZtBoIsSs+obZjh6p/Nm6fmmdoe
NCyp4KgpagMXE6mgRjMZdOEKw1PJ04Y4bfCxRGaJoQpKQNq+hr4T6WToAzlOLAWN
QXV5U2kGC8AGwavSJOsiNVhUT7Z2xQHFZ0HaP2AjIjPzTe+oHoWydQ9/X/VYJRhX
RLMNzbmjJ85WBS5KYfMYfdf40IZDyq700oxuGScItAII9Jikjt2BbMmZQ8UZsDYN
jzVldpbU4P8VaOmOD/ZDMYLqBaqpYcCWeKYgaU5J+rzf5k7bUnJyKOSrTk/qFzGU
lsLzkwkZZMU57vcR7UfFnWXVBhps16s6RolBaD8Mp3FwkBxtD90zKHic5XIx2oQL
LuR+pWP/tTTmCzm9zPMvnIfhRtYI4R11AK9/Gf95jxfTKnpIVWGTMDqrRsCiHirR
rPmVNEEdWwt9Lw/1q5fajXvNUCiAXru6iqySpMBLE3W2tzvhn2oFvQiHH+7QGom9
b38Fr8j6+HxOWS/aqqnmqoB5eQu4TAt0zDfNEhkqIoXqXnrA8DaQJ7KCaXnktK0h
35IZyHiG4ODvf2UjU23VKT4sCRNgoV25+qxACsMMdJLTdvkII5cSBo4GwR9bI3jZ
hFPR8N8x+ooP0u9UhLS37RNVS7ytiR5z/5Xp4ecmznU97n6YpsXs+KIVQp7r6BRI
3VfJmmtT1IVjaAZKXZJSTXuw/fhiFmXJ7VqSf3U3+ZGVc+zOUbdCTMGuQ9iEp3o1
dNKfnIWU/LeRC8Xp6IeizTp/mV2aPJkddRYirWeBftPYpQx/YkRl9dNZzwihVmZy
XJMN3jGHzKFbpqgyy3nAAoImSSI5O+EjNjdGpFK9eWVxI0JCTEP78AzPw7buJSAG
w39lLw3gsP0MpZro2PlBwsFq01aJhIQstpUMx7haIcskqwQF8t5zVxWKQFXW4S8A
vQCW26uQ/aniShmeriGPS90Y+e39VXh6QZJo8HfN5DD/tX+6xbaNHN4KNUnIh/vp
7hmn3ya8wyD1K8L/PbQjwGKUOHiavBCBWxPn+JB09fjvu8VGWu61p4mYf2uRpvXO
IpdbjaWXXZIqwJiZ1tt04EIPlgmTjFMiaQyd7uZpbYu/XjSCkBoSiUrJxW/8mDzz
5aalGs4wo3Z7HgBDuP8OfV/TMb9y6luSFOSRERWPetTHqQreX5xFzdMIJev9JdtP
Ot5OYTWWq19DVeZQJN6I1aC1Tlh+S0FYMAPEkam3XqkRbjoaZnbWU2Ia8jaEwssp
9T34/3Aj7wWCu0+Eo20rjxE2TNCP2igTVdLjqTZ1rM3H/gKVTGRWRs0UxSyED4j7
rfDfFjH/M+56MWnFaLheXXumtWWmBBZLqF/NK9+WDnudAFYbyGlF70NNWZu14p91
5tsVawzRSpM7Mr9PZDbF0Kbi98vUAEPR9ga/QKdUChTvWNz/mxQb5dIh+U4r5w1K
u9/fd47gAJhjjeFaiCbwDQtF5EILgrhC/gN7mR8Pf4yzSeHykT8MSX9XPF9XwmM0
OmanQCxDgFNclRQKqoeAPTBPsCsUHDApNls7q2LM9eb9WI+6vCz4+5i3etJV7DSa
924+8CasWt57X38f3O0jSHl/F9qQEcLXbXdKTxl9IBauptPRiFUDzTGjqsIOGhou
ggcGzaize1qv4U3JE5zjnD6a5XLr6RhvoYWKEopv91Nmc4DBKfKPj4L5TRT6ECfr
klM42YZ+bJTXEq7JY6S4rFUl3UkhBVzukYVW9R3SWk1EqSJzb+BFA+k5itkMEGI1
U/q/CJ5Sc8A6a3pk9lJMpnObzgq/yXPTSNBe21+R8sZlIM/8YrqjyZBWiCrlInfu
g9LOr+1fdAenLrKZryXhtKs1cHhkO0RGv8WKL/fjYbA1lvyx3ivXHa+o/9IDprew
W5AMvrGfcFO7BgBk8uTf218pKyh/KWrFv+5WEtytW43vAMQUo2JCuwFoke+kKM3q
bzIvzIpUPqtp7MttkrklelEnxRUwDEguOpsgiD09dbLlh0g18yf9LK2PjbrGg9yO
FX4RJoZJ0ETNQrB1f0cNd2q4E9/LeOYW/VGFHfwCHcfabUofpMCD6nTXTMQ/uJEa
9tUUttzQcZ4qBiV9V9oZd2f586SrLA26WfegcxyRc9tXiUQ4vpEfiRRypFvRirwP
PJMxlowe2lWBrZ+M8O/NzTPs+C3Nk+TUlhtLqUPhGxW1dDgB3T7aEOcHrSu0hbcM
+Guo0ivewpicHc0Zy95Lp+UD08kMwbbiNthxztf/wepDUfsI+KZ0uCctkrC3nzo3
zRXUGEmDUwri+yUuHe1ogX95OEWgD3Fic8+3k9g63+lhU7O8dknZ0qRUTuQ0Waet
3Xvm4HvS1E+bu5Z2Zwd3E92DBFz9c137PDrck2BpHrA82FlO/m0gw3qbu3Lcclpf
fxAc/QQ95HcaU+b6xD1NmZxNrS9xztjwasVzuLeGlJsHKbeRLY4NgXqBZ9ZYxKnp
PMZzZ6Bg6DAdhq0n6ejycChGLaUd5B8IUhAPxDWzTDyT/EvjyWCinMBgniejo7yw
Nang9A1U/NpY5lZ67SW2zBWNzUYuy/qzv0c0P4sgUQr5pDmeJ8pFXS3zB9eihc0b
HW1CZYik/0uncqOBtoHTxLScFCrAASPYLliQ+UAfCvYtxHUwhZy9H/L4fUwql1UM
UUEYbAxyuPn+0gUeiXWoDgjHqr1KewptXwYDYQFZvjfNgaYIyRfOH38hR0//iM8T
L67a5Xgt0N4LUmX3AlChLVcjQM8sBQVnsNZExcFwnP9SDBgoBzrwxZpWIFR3b0ci
Hxw24tLCmw1tqQYllAF3SIoLV/ptkieNOUvMFxqx5rcMXmgyTuRzE1HR1cd+wUdd
dRg3OgrJSyAZ+XUGgLeHdpkGuql3kQ4mDsg+3yS+nx8Y9hsgglkE/Gz1Qiz2sHPs
d33y9CgZGd9Z7s6NK6bTGfEvxKXVy7EasZTAf63Nkt01ja6e6syj+OB4YfPpEOCO
Cbcm7tmYPaAIBpx22vKwCVBUH3nfh+dVheNkDRwcTwOaJebKRdELElXGSGUKSdHH
7dfIGviKtsOCTBwoxn8M2PX8Ssh5hJWw6co/99NwpDVbpH+QP/dCC6zOnwXjQa5A
RDgbqqa05COWqpfvRRsmQFcAJGZDsd2s78OC3fwUW/HRzFxHhhME3CnMCCTKaGlu
QQIbVLMyz+BAQ+p9USLyTmy4zRbrwmDbfDQSa7PBB5fdOZMVkKE1QH6qlWCeKcqj
paWMSahhjV6+335OnKbAwxLtJhH4spWcKjKWiKA7+sjtq6rFYXvlTOqDTJfqanRT
jbvf0lAf5Tx4yOLrhU0BCv+q64rQRS/J6AdPSSREha1c6oOJ6K+KPWJAryep1OKg
DMhoNso3ECdK28smV+wH9Ti4KB0bpHG6X87260E7BsZY9ai4PYiOrAvZATtiBEeK
ObgbyJKT5uG1n37KxD5m3WCc9ULD2Ki0Q01t5cnwenxdWdESr1JCD+PZ7cnfD5lQ
hFnCalRLAaVJoAuNKteRx096C3MW1fOSuy47OA76h2tyY7ZF7nQ26nWrTVoBBE6B
nWjePFJz8kIoDpUKKiR/WtK3VCKBm/wY+p0+oxFQDqdsgBU+8tHMEwtTiTyyKS99
MS088Kb/owP6uxkaNAcYwvJV6o1OZ28m6p4R+Kn9ndtAyG6J9ggEGkx6tAXb1Jsd
zg7RG79B51x6hnOWyRpIQ1Ixthl05/hV3cy+5roAsmyGs+P38qZn+1hJyZ34W1V+
WrUaQHA81TnpY6uVU/kvmbCBLGY8cVMR0RKmPk464vswpazUSupOq5IHB9rN/AtJ
TAX+aPfA3RnwSc4kp/KmWO37AyjS2AwBByGSIiiUQERduTU+hhdrG/D5Bu9kJrn6
1BEl+m5KcqQDHmNVjaPbGyunsbJ8i+SmLJj00tG1gTFxyxfBXAMrp05xMNtNfFKE
d/vMkKJ7zZa1jJMWG7lcEJSKKWuughdjw54WKXqEsOxeyZVBMorU0eVLnZaq42eZ
17TkcK8QK22LzVqkL4CV5bM+bPqJa6t9XVnvKjbP4sGLXt/gbzJN35S6pTB3TJji
tdi0Il2ys7vfXzoReH7LJUt/6bPmJlYt4gwwYIvBpjl0gRGpZ3Yl/EpZ2Gn17UpR
dfydxl8WTYn4MFV+f44f9jIFNGxQyYa30+QmCnnczVBpajMuQTU/mS/LnhI6oJ6I
JMNip+5KFMuB0zblROhtotECRpz2++ZYaL8A7lUXuxNz2Y4LCFhIaZ/xT6aA+D9y
qTRDjnIOIBLISAsKGFeZYs0UDX33xB4GuQTStpAzWPky6jC3OASV5Hvn5wQWS5bQ
j9YU17OeO+Vt7nmoyS/1uTLzPdn3n7i0eYRPTeSnu9xga7S5pwzfhNusuqJ+QPmr
MVSocCjtR8UsA6+dGVIffeGr/Tb50jEzrF7ZAANZSuP2SQzPbfbLXeGnaOkWJuBi
0E7ZZm8n2+KH0+m7MwP4X673mMgMNBdpSNiPX+hw2AxZS/GxeYOiD3DX1u92ETPh
HtlkeAVqB7t/A4fJSIjWyPivNAWjx0YSg42AxqDxa40hZU+uI/SC/0ihjkVdqCIA
W6ldLxAJYXe8J9H2aVFP71N0Ia6BzvM0R3rSltARboq5gvxnS9zQfN5GM511oLwM
rbdWgO7F6yF/0ISS26vA/7OxpwxLk8RvfT0nxIKEr87DHnPN3D4rWdEW2Ks4dvv/
KYvMPFc747Nia5AhjHGEUlUquJhigRUVJzjgvqEGoPsiC6EqXmv6mGOGYWU8ePZi
v9Dd4aYaF8LvbGNC4phDLPXMbUj2GGk7Hh+aWkYYZaHEywRTWZ89p3NEQnMVgqfq
lkqKlpF+ecqEPTpGuVeUaHHgQ5Jg5nRVEcD6pYOtGfb845gSDJ5saH/2m0LkmaNb
PP07ZwZcssr1SHNLlNMhFBPXaRbOWKESPb3iyT6N++C49P1zfxVlJTmbLM9MDQRG
9jjMsJg0oiAUalfZAqHNvkJ+13rEJlmf/llULXDoLVXbzOhCQjJdsqA4HRMaaFOu
bmEDxUxHL5Brcl0bdVl5UTdnVN4abTwFisHk1atuuEr1HodudM8Qs53nRlf7CMfj
0BrYR1KOxsR1b7f+WYpLIbcKVFiWof431RCv4MUsFKlAbHXrebkFfJSI6OikbagR
g9pQMMTMCDGkEGu+HtbDRJF/iHkwdTM3FpyFmPauFBjN2s5dYBy/IqtKJmRnq1gQ
g4Bbx3TbuJZvEN3Q647mZLJ131o1DSMoMP/deIsiQYZ4Spq/kU1LUVCUD+SSHwwV
bnR/eBQc0MDF2qj20v4guIti/EHQciViUN+C8tSggJypAWTmHtzvvGMos0HzKB94
RKvFf86+DayLfuKB/rT5RT1I9ob7ckXCgjFj2aQr9q+iEnz/WUf4YHfdLdDxmmbH
T/JFHQ+Sas4yTxs4IKECSfoOvvRYQeObM35np9pwTwOjELiCJ3AvbWnV/3Oc09fK
NpSOr7Ko31p7CKLMu8n7so2QnhCXLHtKrzNI3GVCDrh/jvqUtDbhsB/87FogIpo8
tP87Co6bPH4X3tPW30GlF6uGVZboDq+yUsc9H/UejQyGUD+qqRlNq6y+dgJMHi46
VWksrtlX44XcF7YwjwNvr/WigZ+kSQfnbj2U5ybfnZJ0+3hrenIBSD4LkNDpD9d6
xD0iY2jJNqz1BftcN0eV1aNVXQPMX+tRPhS6N3rFHeJe9zExUTqAaeKV/uQe+PSi
7uX5C4t/skPv/Wzt8/UpjMSSvPCsNQr0WPwFXL2rP7zNiDl9u1+jRn5QHYwsQv4H
6sq9l24N6mRgDkSy0/r6+Zj5KPCC5mRyH1I/0l9jrBucObano8FNRS3IJaH+8oPi
VK3NFCFHBnaU4gbdSkEI6UMvp5o4b3VuI2Yg2KleV1GYtcKDgCyi6x7E3VLByl0E
mfWFCoh7QKX/rBK9CNRrIIkMwINiLaBZ9+B6d1y9CKqU/1jMmmMoBoCoiEtUhrGT
qW/dP/fZA5sSvGW6wPLG3lB8SNYikNWPtEIc7rX+rDN/Ynt9YGCE7uaum4Sg2vbh
RXByALZ2OdYrS1slVcZwEDB1rBIPnE7urZPs7lfUxSXaXEGHe+BX2smMgZ4RCHZC
tUBCH7w/4cB6IfzTZyY9qzZzJ+V3kRAG7jVmh3iWg1yZXXZFZGEyA8XxYiUCO8Qm
by39jCUDZ1UcehIPpWOYJiiA64DpArh6vxmjGPYIewwZUxL0S1IWUD44DHSfJoOW
AsrQbicMp6EF3xd45mrMah7qsZEy0usJteszZJVmY2Qg7+4rTejFQ9nRDBVp1rUy
Vq7HsvCILAs3ZEAsZ34SOZMWrr449BhSbuPQRZaVIKdteg740OyVfgDoa2uHRGRF
UgJY6gdgWTncxuH6CYD6AzM/f/sPwE1QXVQwsLsrFMDuiGDeB+NTbzfGb8mmotUf
tm/n4eVBo/kdzpvYa5iGqZWERrHMUzJFbVQ5mPzgC/LSZ0+emNLXoCNvv6O7QJfD
uIrU9+tGgdVaHnd4N9pRdi7A5/A8TkqA2AfItSSNKfQtkSJ9AZpYiKtlKVc8pJ+e
uRSxCMPzIbeNeIRu4oMZ3AbIwYZomQOcLPyMu5e01JlTjkCz/u3aXwue9t5ei8E6
/TYxaGPCBwFSRQDZvBN6XyGGHTFFZFMBrN+VrvCNYBYgxtl15Ft4d7g4nC7c5OP8
z36RzHplM23Znvc//+codzReKZEpu1WOJgSg50rnRbVIBaGt4mbTz232HKQ78ClL
GJh6/kvzxT1GOBsVBdXuH+EGSJVcjl9J4SrBeWXCkBTqd+X79P5VrKD8xm9UxuKo
aGYSafLbBDJo9flGQtlL3iP0K3Gfa8eG7GsE65bjx6JkSpffwrX7Plk8tZ86HJ17
u8xKZQix1ma0QNNrJyvM1Iqt2Fe+ccr5G8Jq/nFpXhpyY48yEU5JRr6rGvSv5iWE
af23kOPUvbC3HhOYPpb5x0JRGZeYjEtNlp21myVfywdFSIFHjHAqlxaX6hzVRiwH
gY9BDt9khnwq3tcv9niA/xU5ZY3kVvYWchrcvBiuy4UtQt917X2NiLP0jrThjDHO
eg3V3bUKLkggdIta+dLrh5TDdJfxkxUCaJttzVt/6Vs4wQ4Q7k1aT2cxOatzP09P
Y4xCnzIIX7uAlMZB7Dl24ku4c19NbXXclUddvzLP3Ojqr3smRrL93AzaxKcPYdPz
mPyQ3KZ73S/QqRo0UdhKn8Fu9deU8oIzjHMdTbieUFblNCtGvnVIUOoTNgh2ALmm
kALXDViZdu5oaOY8OQT/IK+R5jVIrqaaeo6tv0UtWpMknwLQ3vcl61FBO4RLqnT1
joEOxfcvzAPZ56H8vf9eKehBZTEfLqaaZdSReRuxfaZDozXnKYqffNz76vZ9D0u6
xAKi+zIw2/oeJg+yIWWT16qpTqxVXmeE6cxfpP7Yl+IohrZZ5AytafgKPpHBbBir
+Qt8XMg1A9ZpZxGShLsntlFdxyPHSUY0nDv3RzKsrrk2FSG/BwEM+TSCKaIYjU16
84xtEUZj6RFQ9JTvHg5WbLiL43X851rmjt9SDJBULEGdbsMe22LhmNkgNWAAAzgc
fXenPk5Le69awH8lG42jsPvZ6aShHS96OXECXkAS6HPx/dAakS23L4vRyyWUJtKA
FnC5dIwADl/8nCN/jQX2RzPmxRngkWzyBbj7RW8ryYpDV1E/22MV7ipZLXoJtgwh
Z/xOsnduXdXLSjtBrChR1uZDv4g7P4Am8S4VCAYWedeVNDgfkuFWTfK2vOkKfwMK
Tjpgkza28HEFcKSd8S4hAs+5zRR+OFw7D1F3yrp7LGTIXv3cQHd6NlrckMQMovw+
IcathK9oG3xJEW92BczP+zio0AGHHyjTO2Z/twrFL79xA1JDEPJqcR82PMciwATr
XpLDooSnfssnM2f6XfJXSPQDQx/9AX0m+cUT7D2BsoLB17EtcWv3yGrWdfzH4UCQ
iArnTOiZHc8hKZI9lZECxMGsLb1hULb+/yZQ6DJNTb48XVOzz+/PijWibjghEa4N
qafIxF36xLrVcPdVFCjLJnRX9oDHrFBHwk/HhpwJ7zI91lA0QY2XMAbQJpwIWtGS
wGSLHC3RiOuFYlcAFp0Q4hWm/wEu8dWrUZDNoGiT4Wi4eDpQluAL2VRXV5gR9WI4
JpclEBNw/FPq85Cl516m6C35HRJg5F+VOg6xD0fEqL5O2p2BuJ2h3c8IZWoS9sNQ
binMYWVcreJhYxSsEvTRVym2FyWwYX7XEEmsXzKk7xJrHAF72ncgYuPplIBp0Sdp
q6P+0TOQpWwU79X2Sc5yybet8sRogo1rsVpGfnqmKjyfskwlYmJ7NDDHLKhEiFFE
fnBpGequotnsXpXLbEeQ4bkYELR7q4NgXviltFzdHJxLizM8pJ+hd+r48DsOnOvh
9iVCKmBqZ+IOUlIBErE77NKtjWS+iReTuuFsDCZj6wLvwXV8kxOyeYkhvooByJx8
N21PLt1ftzLveTedwogh7UN4dOLnYPzOzW9rXjtSWKeK/MU93YfGiSfRxHnvxClg
kjODX1lADm9m73mS+aejZwhYFoUUQeU/q/XQW1vqEZ1s+gzdIh3m0FFZENNyw72P
nheresHyHDOkjTm3U7eGaJ+MWFbfTom82a3gO5/sW8aCOzVwtFSYH7y3gxwulNO+
lXw+HALTefkgftYY0mB5cqIDE8Dc+/Ao0vhlPciz5Lksm3eg6/S/sgd2XzsKBvTr
5S3C+SpzwFSr+8+BHYaD7TGiPfwoVK3D7FPoO0WNyGSBBTXSPWcAvWIZzwzuCDKk
YpAz5hQosMKdlGDpgiSafnK7DFA6elsyguTP8gAhAkWU9jiA8YeWZN/kK7JH0TQk
S09zl4HhpQhf34rkwBk4ltJLglCsqBK8fqhriYcCb9O+tHX/eNYPt8NZk4J68zoo
xvhRxbCxJjAPS6B7tA42uQ1gFWMevFFMuPiHXT0fyM5CnDIvnBEFjyGZ5FDh8QPF
mTKy6OCGmXamYPypQINJB5vLjms0JS/Ai+MxyKEsCJrECsWOD4BfvMybuR+QHOal
m9vGHtx+wvaxBbery5aMh47wMCMPooxnAErlJEXh5hfHSkvxKatUg/ZfahVx7thP
p63Zm8VSBeXfDZmdUkCq5yqnt51TXk0BTVvU+MXjO4ryOjkwj1Y5/XitL3gZSome
xxkHJ7po4ilf+T+rQu6mBwFXGPhKkXdNp2lg+lKePR/wgb906t2uWj67r+nvhLuQ
JhTWkW/EdBvUf6bnwDodR8dB9IXv3HdbJ/OR4GnsqBFQN8Y/x8quIKaFuhlCmQ9U
WLpAxwUzuW6ZivFufqon+wLUs+GrynJTjIjxPv38FF3cx9aOpIHJqd9fff3/Hd+b
pAgJo/PhI3XEInmQr1/H8pnnG6qOi6/F5IsvwU9QTwdemN9Px5QJ+h0t0rPXE58W
4HGCofM1bQCNZa0ry8XzJTC7SzGlv+3VUAib9bgKPdPcJ+rajQGVZC3Dy7n+ZBQF
9J6rig5YrMekBvN1pCML013ymtrCOC8Pqx5hwDgtIwkCf2twkflisMwSs7sXysho
o6MLksXO+3dD1qM8RmSywYE/Ump06xJfzQSFc0sVeg5tXexGv66u0ZyJkdjmfdgJ
+UCGEPjdL5ZSwpgZbH6tyRy60IWxtCGvbxzWY+F/ZFKijyj6AEyEmeRtssycrMev
w4qP+f//3EMAPUDQOE6n9ntPMAnUHQVv9jb4AdueGdl7acnc1Iusih2sepMxAbNe
JfWUoKaArp9ov/4usCo9kq4ZAKIvcl9Vmrd0PIWO2yFKM3MrgVDqcrM6vVhCvMc0
l/2N0RmmVYidjpmTdoZ0UaR6UFhC0bM4oUw9XR+MabahDIHcM+7a3oRXUNkgWcL3
bUf9GKnDzjhs8uVNLu7wR4oRMadc1ntPiK6bL9kh8VxBlT2QsPYycASWRxiNUrFG
sIZDDpEasKVam1nPMZsXU1wJox4c9Jw/sgGwRuctBlXPDxLrukhcF+T2r/xOifOL
fpRlt/iE2CnkatNg1u/xehzFIxdMC8f4l3XwjxhYsYPhWX9AlBp1HmzAksrxeV+l
wpa3hv7LrVezWiC6PBdM62kYWQtGvHPYAqOcrczDoeJd4VmDGbiKG0jaRflk0/N1
T3jOgP3nueJkO1weZRk4aouQabDcMfz8qEGKRFVI93pAHcBxdcVKzN8hpgeWg8aP
4Htp2Zp5Ijx8ZlI1S8kHS7xY3g6EC4MoTxH30u1fuYfJKbR3/cqooXwplGiZxh2/
YNhU1SBwBEcKDH8vxtL1Jt0imjCuwlAKPTg8JxXJEjCbdcwAQZzeTtMe/JHsUi/L
qpaL35z5fVtWco73B8od/2fkyMkWj6TUeu2Xf1ZgSYfu9Rr+CcCXExZ+DO692Imo
jIEqrjePSRni4f03YRo2Vjri/5XFGSx9VpVv/rEW0kc7HYpjOSOCHP09yPYyn908
NwE5CPGNBhZZi8WchYvU+TUez5gn0ofMWQrzAfn/5ANxPvN7IKOWkeF1Pskiid6n
TUUe+7cdDf3iR+Y9AxdbM0j3M/RuYYF0emlfRPKc+VCKvK5DHy3w3tBsKSEnsitW
DREISC03zh3hV67Kxv6sFTR9A+BngAKKWkhdtqUfI3DH+j3rtn6oITmn/ZjGwTQ4
KUWEfpbRDNV7CufHiQ00UtHlxQ8RLSiviGwCAEmnqwz25CsUsG0zk6dcSqg0LywR
74RBIw0vyIofFQzL5Hrgt5wt4XVQUcx24b6ixWUrA1LP+wlV8b+EWl2GU56lg/Ze
DX+Th9127mzfwlF1dbEgTjxonUsndoLkp3IP2Og/f57CoLJttQeCdrwbEXKl3k6v
+9qd5zImZiQ8WAyRTwYFJRXAnSFlPoGVEjvk1DSlfZqaneeTSTr9PyUW89L47Ktm
QzaScI5e30oSZqDnhKdIdyH7eEJ8iKVn22TRK2Kyq3of4ij7YgNWd+G6A+rrIuyy
V50VRJKOxm1L1K1XutysAdcyAikT7wrsj1+H0Ds8K3Dd0LQlZYpyum17oxxwnOZa
ZQtCPKiNmsPtLrP8and6/J1xX1yf0h6dqOpdxRP20E2ymJNoNAmLXLeYjvkCij0E
SSThr2mZBy1sqTNr0YbB/zsQkt6BngcInTIwhXcqAVW9VJuo10Gkl3HF6APA/c6A
y6whvkAcBk3nneb6xg9anU13MTKMoiy6T75FUkIQsrF5GcrN2cuG9WYWstcPeZH1
oGFD19sOqp0KAwl3meLsPmTgiHwijf99UX7Y+Si/vN4aHy6nZrfIYyAJ6x0nTFaR
4b3xnPOtjDDjcu6JILt4LyGm1Ihh6pwk9PyosL1gAsWt6wJ9CC+kPXcsCp6/6PsC
KzIjXPBb4XRmaODMvqYu2+NAO27Ay8G9hgL4oyfO63FVZqFGAFY4ZdzR7BpPB8dD
a9CGk9TMWWYxjaJeWESau0nOhVLZGvaIbMKksXs0tsDHIW1/t3V+0TWXQnW+xEC/
SMSMlclvToEGIJLMDxSuMrLTBaxVqqHFZ+QfLUYNBSxzWCAd+6RyoDOydpxDGgnq
cXax/222r2tybHbBlekl7RaAyBDVjzgnaubA15SZMv17pxHj1Oc7Zv3GWzHrtp7s
T3OS7SHTDLxFfnYgKN6jSpWRKCIdeG1E30aaMGmD88Wzx0/DkBw48+A+eipumg7s
cEwEP2xUtbYXpBr3NUd/Q8RyJ08S/i92HWYxckWMZmM2RwBbU1cuNrSa2bgwaDJY
UxyxBNTBq+cnbfOtER6h4UwJk+D5kPJlv7eYDGlGD1qqLQgPysA5FIYrvMHwb94W
FzJzk0y3CkH/og4j3ZtwQciwuiEj56j5zLtKFtC7Bd1L73FyRK2h/eQHfVKx+aPJ
cKsKdeq0QaaeYhxn5Dd3OCHOU65Ksq/U6mv9bszqcF4WsFp8dz+XFbqYQRffRv2J
mbN2xEmOqYlW6LTnyqmtCdfyKcx+AQvUX7zGa3SlsHrjnEfA0aekWTj83GEA+v4+
awwMqhLdtri9RmKEb4rAGvTlOpE91QGJCjYXjgLIjPwVSathXreqHIwovGHha4vZ
/KCfygzG8IspA8Y3uQU4UDQ4nu5vtjelwoZdG3gXMwQ26kHWI0E+0xFwpA9M+ztS
Ro9NSSHlPp0canMebEl0tPx3ahJ7XLSDdFirTm26JtVjf2wuJ/Q4l6XKb+L1XNMy
ddCQZzv0HHKUu0tO+DVtmvlBQ2A/ttirWkwxi1Axco8NZ9bhxqEcr/2eyA3MjW+p
tL9Yn9rvoMoTHXtyrysbL2U5jEQNrYpF/r5GAbACEo02FTS6S2qUzhtfMkQCtc+p
flqQqunmm4VKzDoox5DKpTTb0LsQXi23O8fTA18Kuhu4lqLaBLcOwAsUcIhlSO0F
ZcOwEHK64vO391Wg89tMw+wJ2wZMKaTYdB1nW2GEBy2+/5XEx4Oq0+ZaFyxk/s2F
Ihrskph5ypBSDrw/4G+pSMAf9uUiLYcXfdVUvGFFv6768JgclYOb1nDKugAY5Xy0
2AiHW0cZOkLBfMvRdI2tblh2GI3ETbiXhLZ0NaBv04ny3sXbZhfu1aO0wckGhnbo
LouBDOZL9pRy0HOSuGT7InG2bpUO1KEeGLo8vTxKvIrP4OPHTO1FZepRvclAEz3i
sjpuvlaspNuB0VtqEMLyx+f925VKTTmfBeA1WJltb3KJy5P6V+OuHVi564ag2M6Z
d0xRGFqZMpwkh06LVhxE1FlV6vnCDDEy/96ZrZjGX2K2k7otRm2e+U7+xKP5agwF
8xboY08Y7IBWCZb+moWZwnGUJBSswg3n0ZGKtfLKRHYrlN+fB7u9uNPhrJ8iFU+j
OdFB1oPP7e/T6nIQqhNRHnWw83DKB+sQo0Q7ZYGZhDWgW9y42ICaXFSgkx2kBopf
L6LR2esS/v9BSbvVNwkfXBchgrYDT8hpFFN7nr6t2GipOIWKK/oDTePF5NdCjOC0
l4QSOgU/0I5xxDP7CBnfDR8z4AJCYjosItn4btbizVN9OiFKmiN7b4i2aQCLZ6YU
1TfbcNmKUaj+y9/eoqKG1A/1uBnDxs678v/aw/YjZylAHAQmgc3GR3kSSLxoAm0D
w2VOYOdOuphvIYE5ZkjmzTVoSI/y4w3XvuiSS2STo0aZ7gHYhp4ZyBumoV9zm7EJ
FitwuyImRPg6AQm/FY0hdpjoXoHD187ebVDflIcPmIAp0HLWrfK6dCgHZuvAwUFP
Arh1C0Rcb7c+PwcGFSOBJK6z/a0ExR0LcoaLMHr/wbqeiCKEwbdXxXpaozzpDSRe
s/4HN3OF9wEaXfFlsjhOYHc9Alh7pz6qNt1f2MsmxZf7ocoPJ+eT2yUgU/LdnW1J
57VJWMdURVgNWdnLXt6IkPadMZeuJjQDvVI8LMd5Exmvr34p5X3ZuLe+BoPXP+bk
MC8HKIrENSoXsthmmZKZWA+o5OEyba/MZJiwsXgnuHeeGm+kuG1DUfSP8yW+ILuG
QFD+4RMdKQcs/8Po8mptvPh+42xLsNiN+CH9oBGEJ6V1d4QWazm8UdVvBXNWXiRy
yFJWuF2ADgixpT0PF0l+Tt0e8CQrAbuAxbPSpE4TwpHfB61Ykgs+5aLaD4yUs4tk
JnFHgc3ebp37cY++ijzjjDpFeYH2OTBfstEMFYlBzsLRtVDQ3/3HeTXuyd1iL70K
ACutW6OQkSZZhUb2zXQ7bKODkuJG9zweQqExu6tkOhZ3+o7QUOxKhFOlBltSd704
BoPL+Umm8A7YRyB1SOrtK6xOdEKaQ7EmwsAHK4qfcU06kUvyBMIhpO8juoMBMyE1
V8pg0gQa0jY0V03tslTsiDzcQYjo/dysUWTebw+eMQgQzwk67T26xV7fpYZtfw4h
B5bWkPmDSr7YEm4Q8abOrd6LwcpueokZTfkK5vhrCEM5BwTGK04TezyRhIrYdwnL
Ykbgeg4lbveo/RuCkZ6uJLMav41A7OB+HfOIoCbMEAhJj1C92LQZ4PC6IBv/1UAU
gA3u1c6cVm5Pcdo9vQaY+ib8c1751TAzqx60Rw98xgeMuGqddB8Q3NZbv1gzvBgb
KZGixqAXu831BC2vl+k01LdOHEhlrKIG6cSVBnebeWp4PlcEVXZYKxdlqyLHLtzr
+e1kyfOnyVBp7EoR5knUsVc+vUn9p2B4X0lzBrlWXF2vHpIDLg26tPzhtKO8EXWm
BSm869U1zSYS3UkRC/qMaEJX7TX9jJ7eP031zPjy3LNUykQitQc/X7vwAF1WPawm
oC1Nb3N661Uki/+znbPx8PEpetf69phP3Ik9kfLInwu4E6ATMSGC51mq2SaKLfmM
H7nFJW6q5vgIExrAf1PVqB0TWWnX/Cj95i3OoyVljtIRCUU+eoFnrWBQ5JFS72bM
ORRxwDzPd2ekzUww/1k+IWphsmX/ydTPpi1Mo5kzAt3UgCUGBP44g0H7+Et3DDHv
CInzNIUyDqqATwhfnHEkjEpaTqqGlTHN9Bgw51hAR4xa6GB4kTP+8VB7y+7hg8Tk
tdrgA7yU+L2slvPJPzTkuLTZXggLCwqp3FhfRic2vx9vddJNzgLue9FbFSOq80uA
hfJTmlgbXrA97W2MtbhzzVlG83Z88BBC4/VNG8BCigrThqjT+i+lCPptnO+M3sSX
Boe8oWXfOuM+Hiuu0cfDRTODlWMmn7DO9+z1TuCFCqOvRNj+pbY9tTY6hB5GX28v
BT4RdvCPwUxcCvYcZ5g3wCSeJIGQEzIyitmoUqsMUTVbEcbQ55b/eoeUFNW8RLdg
dKj4FpyIqp5fuXvM7QnjE5/2RfOTFSjeatvHIBmusQSdoWeE0zZbPAfQ0Z0D1zKW
sMTcHL39YfjQrDO286jMb4FRJ7CsHGA5xbUT2KtTeXatgSJRT4XytB7W91wQS2qk
ymWhAWm3fnFk2V+QqW+UDlp3Ylhu6+1O5oKoNuvwVVLuJy9D2jESw4bjarARshzx
COgmfkT91MNs40c6AHRP2t3wXxaF2183XvpX4DHTlENw3JiG6PlAbfHlEz1/YeSf
frzvtSy/jdUvnyYWQZe8F6CSF7GN/2pRL6o6axyiW3+WET91IVAaYKnSZtB1jL7O
mZYakwkddcOB6Jlwdn8ygGrGsTKmfVLtzIdBM8S49nklF36fREL2akPN0yOxOnZ0
/EHfSMaWXCtuC7og3WrZ3fnCMbqUw5AEEEJsXeNwOajhju91wtfypB4SNuZeYG/s
QqOkgQQ356TB3wYiE0cP2XSUbZ5e9M8ysR8tfmUeKrZIF6z0TjzmWUGx3jn7KoOr
wJhqO1iqYUjLJGOU52Afrva4eLv0qvnoqTlRFiYSXVwSYVGdE6GGdTrmdYmeVMzm
HJTjkQ8C61BHDEeueEQ/g3cGrnAj7z1/Ob/aGB0u5OwcuF191si6xub/aajVowEN
QugcTZmwL5W6h/n1jo4Ws7wmAB9rROyhlaMKInMFfqQz5SYgTD6UDRT0knG+oM2p
RjhKIVTPSXxPExP47THe7isfUh/i7iyedJH4vGfqNqtKZPdIqRx1ur7lNNdFOcxM
fCrBfRDkoxhRAOXmY3GiaB7U2rbpC2IulO4TVef1xJr/0byT10UxDjdHnhprNjqe
AgJb66Zao12oIP+a4KSJjnhYidJGW2sLZRjtnHq+9Oy7QmB8BGF1GY/qMW9F9ZDo
z7XdERAx7jKnfHGQrvkSOHU1bSMSkcErHULsxXsa3t46Quv8CtzsSBXBptGEIbpf
mpE6pBI1IfwsaFlKeVEkiBPQObPU8bH87vhf1r0GGeame4LSmexl2GiiMEkjJZYd
bnWoXwXfgblppq2mRaHIviW3Hnn13ptf1iNQH6KpY+SReohDV7kZeQw7KBAiafyu
jhl+SOEJ/BWkbEeTjhphaYqoDLwCCbb2gSlea9tP2iKyWcNRz3xFIqleCBNl3hSA
iw9kp+SECMGMc5UHn2KEuw0/KTvplyxzXPHY1LE7D1rY1LC0UOrUYFGFQ/lk9DLy
u8O1IcWNLNsY5hITbgrA9K0wqT88sCWH5Hd+qcs7ZYhvBdRCmVWFXJsRp/mp8n+b
9IL3S7G1VAWeHPuGsyNOVQVp4eEEYMkkEy841V9NpPFIpQHWWinX8ij/m3/yDVsB
e020BE1QLyQ1lVOkXneVl8wAowroWK/WjUgMFTmp3Mnd+1AyjEl4ZSAVKiVEwFUr
5dCIQzIlxl5qnT+QVo3PsO+Q1XQheW8ZEklCHzwx5LCIWemp9qMczzYII/7YX+kx
jkJ8iYkh1rUYoiyjv/unaC5L4dkoZwM1c/DMKcJxqGMs7AJG3POunU9xGa5LxUZ8
z0HjkVpeOnfJ+UWFghsi6yPvKnvXPouuXHg2AhnnKdYxvTa0bVQNpovWZrRoQpOE
/MzHmDjAuFsAwuRB063IUZLA5LWHKvOYcwOpBDfYfhW3vvrftpxojHbiwb0SUTLs
mepbrCutHoo/BtvxGa0+fyRu+aFqXIV9kRYSiIPvHKR2ogtGvPLj9PgIG7bzs8eF
io/mcqLU4v0TbTkxHoNU0JAWa2uhTNsHrY3m9QxzA6Mx7wIcRrLRv6Mul7Hxdv1g
mVn//BLjjJoTikV1uDcuLJoIWteGbeVAVaSdW6WO3KAgipwU3+EB9T76KDSM9Hwa
y981NG9JKR+nJlt9+et5ieYFlMFktRUA6J0wXnkMmFeANtKG1yzgEGQQBM8Dhocw
fnStuiIcb9UWtp/30ic+X787bJThSlksJmcyj93bHHL1KWPlDDjmkbIno1vpWbC+
oVnlFgIqreXcXsGxHmWXgm96GpZDOmUnbxJoVF74eIg36hVhsemLUre4RBvQ7z7U
vQt9mxTHqHeUpF38clYZ+oU1Xwx2e29zJs4MmkD9R33w8quCWagLsmva5a4dXjdw
nLi+G8whzPCX+f+geBTlMMyFZ3NWZHSnLJ95q5WXsmhHpD8U5qvj3juKvco9wtW8
goku6AaP0+bM+3PfHgcKXh5oRXZ8oalRHH+w6FrEQlqXhzffEyOvJmiGNg598EvQ
ntdWljaUKhY0C0R1Pa27LaWZeyLDURGsFrKuA85ZbDY+7fgaq0xIHkSlWdY8C4IC
hzcC6PNELA+EmXCHXgK52zMvDbpJKNRqq2saIkTHq1jsHHvFGCkGuc0UPjxCf/TG
rzO+NyMQSJ2AuKoHVa1W49O0k81lhvfIrFDAKvwcZ4oMPnpW2FvJKtGQZG9NIjH4
0aME7sXbFyv3XTph94rXFnfnJzbiTS9Ly1A/2gFnKUlYqA7tIn7Dpo8PbqRJ9mbp
6ndD4siQUURIy+N7+KvV3+PhIVpDpe5LRCAFMiyq2guM7gFEzXNv6QEadsHcN/LL
wKzRpITobfUctPV5fc1rzNFYMqwi1LGJW/vNOhRUegGnoje+/BloCFUZKdbvFJ39
NIFrrSHdZtcCIXzgtRb+sY6l0Vi+CspYOTVIWOr2JPJATZASJKv+Vv4u30QQ4qej
viswahkb+Qp6NDyMV/5+ZTzcDpEMjgbUIbK5hKMyf7v+RFPjlu+CF0mEbtTj+5c2
CXqaA6Ib4auqpxhsTyz2v+N2FHOjLFQPG8Axp76zY/bVIc/yBOx+/JhimeutZh6W
q3X1Vy+slIIG1ydwogSKYC/i4LXjQmF/r9/jcdSnzJJNkoZTQAjq54e7nYFELA3C
8GsJHFeMdwPprPZiQpqBTC3cGp+zn8MZdK5na7YN2776ioLjRZRJHpQW4fX6lB+r
oYEztFKvd+GMW4LMU93KSDhT8Qm32yjFbwaa8GeMdRTRC1vPpZ0AirIYuzRnzuvV
ATaB3F/fMQu71QDcyGJF6qWuTbIg1rh2jPDo0qP/nJhUHInGM4llNmkzLu6IQY5W
ixcvmzSjaOezisqfC3fN+PzLZoSCDMN+FcFq4GjtzQi4CmXmM/h9MraSxy9+/WtO
Yti9QA+sbgr430kCIFQxJkQJqnk98f4MdJ3Mq2THQF7ukk3/zF1amlukYZj7uuz5
5hHHRaQpnc2Hiwj21y4/R6AUQ/lLUyXCO00cI0VCxjGk97pdGIkLziV40NMAEeIi
tAgxeqDWiXTHzj1dsUJ7wJk4y44LpfS/GdAMugjoKzesMxg9luc7VKF8X6i9d6Ka
IA7H1L7ds6rJMjlZnhDLrgCVIvoIkhfejiK3SDVH0zjkAovP4pFvoXChgcwqfYDc
VdINv57Ml0fDlME9Act1/8iH2ncEg3k4OggHI1UTfTEsuJLV18t9HAFGbvm8nm4j
BfzTatXkrkqUuIGGMxAcIfBUvqAm54IJQ1w95PUmVtYa1m8FG9M68N0Rsx9WiHcq
SiD90h120IWBe9/3QbigDAsy4JGLNQ4wQbzPMQg7hUUFCzhOCxaMX2RILP/X8jKr
7+iyL81n4Kv412Jw1g4Pswc+AQY5R8/tAC6NBgkfISpzxJLahxdcYueqEXW0InI+
HkKSiZjqXzAPlyK6kKU6X2RwPmIvf6cM4Z+1OXCptIKGpOkNkRLleq5Ens4ENVhm
j4LZKJuqK0JQNnvTpBk2W4y6vw0GsSW48bTxJLKU4RhUSQO13uo5jvXOaXseQ6+c
qVvGx6Wy7h81srmRTqnyAunBiSw8A7LqFjQrZdvu4ldLsEJmFQIRe/njk2QbtHxb
A+OUBvES2hFZWe93iH95o8oVzIU0Z21FjWtqqTV6EdwjTjeqgVwUE7/yvOTo045I
HLQY/0iRhFZ+7vJl674dQqNyTiUjvq26lw6lZqh3GjEZKcJRto0UGs+vNMS6+COd
VHU6Ssje1BBdkFU2i/WN9UUkDbQ8BDyBcuR91smVFUPGv1xU49d1C4abVPmUT79w
jY23MNRZUnjSZsIgNlrW05ZDAsKWR7TF3jCbvvmVq/EdyYKCwZ9YEyW4yljT3pWa
jMyv6rqdwWsVXJbNFCqCRSKLieYHlWdUE9Zo0+jmNAuPDu5BcF7n1wYUlzNoSI8b
+5dn7hc/mNViQLeiYwzg6iE0/XdLQu9khG2Ntdosmp/bSLztZZwlMibKQxpDtPkU
69CZUhH+OB9Y8G14GkiZ2WEWnpw1jO55BhOHtRfpYnHghbQj+OO/FvaLhxKZReSD
cp3HsoqqxxV0RFWdsbtEQwzPHWKIVOh2uaPwPHVnj6oFO8SP8nkgk32Hl3/HRIm4
WFddYRbWn5g/kiOvhiA7E5b/v/25AAE1NRKQHh8lVjzvAJMHs6Amatp0L4QVEtfZ
vTMmW1mMbuRZIyhLFsRSMjBSTLJExN5g+r5yTQworcCBNYyeLZL15jfJ/YrTRZ3X
r2vDvn1Jmm0Eadc3Y6Op7E+Sj7k9HqB/I8bkqJ4VavgBBqNsL1Dgfk884DduPq5N
m5w2Hu63nAN6cQllOUHabYgcyEvD2xdyz1wO26XGJOJ5cjupofhBgCz9AeUQvI1K
AlpuuPn24dsDyVLLMxTxZh2b2MMpm/t2DKfRW/Xst76gYMxVgrXO62yZBRqNFaoV
gLZlxXS/AKmED2pl7wbM0zAqDG9YCqvH0Kk/+YxG7rqecBbCsHl8sbR9e3uTC1Wl
YVKeWfmYjQnxvXfsUG/tfTU0TPGYmlHX/T/gILxAgAQOpwh9g92/Ew3hYSLwpSHb
ArHpbVXmb5+Se3rPezGxX04zeVeqTQjGrbEKr7O5Ivdwa2w2PP5Hn/TxzLKEV/AX
mUSBPZ6oshvVRW/NHNfB839pf122z0wI+/tJX8ug9k1Y6UD9vBaWPtkluV/QxgBq
FGPZdpMDqor5Etw2ulxhLBgejb9QSIuLUIGHtqo/eHMZwVvYjWrRYBUemVYzuxvx
0pc8WTbQ3EwhTml3JyuI9DZ2AmZMsDaaXX3lnPMEFL3zFSS1lbEjZCCZEs9W2FTt
nrG5QaRezEZMixcL6cH/Wn5MLbzAsbBRVNXvKu/dQHnI06rbAwOm504mXd+GI7j/
bK8UmnDVh9zP6B7Ef3T5EyeolN91c06COJO98K+T1TPmlI5P6gPsxG+K3ZzTGQ15
ImmBKzQN5Of9CyhFBg2rO8TbEG1vtbEUssq7vkc7fJSrjE8JmjsyUyYkoOdLkwCF
1v2R8cR/KFpPlz8v1s0vX9KIOHDRrwKn4kfTuGlyGHEImmuKVtu45UsvjeJVWg/v
efESatyiH6YT7CSWeyAe+m+4LCxmJFU7ebTovVkmb2zjyVqKfTSB3HaLE9dLi2D/
5RVOncquOWFtQdK0ZwTzH6LpM23FyzZZYeFblWX+p3FIJJmXEECGaXMzCax9A0we
wMRfcXiSrwX75YrIWMYOKJl8cUh07nOK4jEre9hys57xFOSl1WTU6ciCre9weiUJ
om0U+f4d1kPF450kic10E11LybYjbJDuF/iT9rl/+lvPbUnatC4CQAIpd/Qz4uRz
fGZr6fGB+MD+kl58GOckeZG4qAVrdvBduKIf2qpeJ/SiGAsmTdBrlMXZ77mrr/sd
u8LNHGOQwJIN5PZ4GkpqluvM3S1JtLiP+Cp5zEFMqUUtgdshH5jvExLprJxyEbal
3sMyjP8tsJQub06Ih0Hi0n8fjNmtXvvn2wWgeLsuJuGSq+iIEB5QLfzh7WNxzpxX
NBWIDvQqTlDLYac7kWiI5QIcdlPTOYHsWU5LY4BAhCI1sQCAOVBTDG3d54cwp2DV
/8N2Piv1rM8cSVltI2th7iXDNO3BwAYhPPzsLKGNkqGCp3AXVmFU1b1K5LK6v+Yq
eFVteZm/m75unAAKAfF42Li12HPl6W9DsHTLNPR9fo8b1MYnt6RXbsGku01Jfpmg
FqWNt6Q/r1BOKuIzUACNWXiagEj7pI0+8zkmIokJ65IvDGBb0C1xEr+4rq3NlxdC
jMEdHjyStJGXfIyNZNGL9Xjoh+Zf4s4bGzKNgMmc/gZygjm2CbSMByyC7wtab/xG
8CCH5iSSxndYfCrUVOXkjUDxSjeSAPWFV5wr71rVIrAn4x3+M1VC3fl4CeIdZDjn
WSluWyI72RMlwS+oEW9sqJW9f2DcaSo8ERl0WPL8iy6pGXR6Er1bRei12nAc7d8m
Bf8GdmWOYc29uKodRY5LGPuduv3ffXZt1t3BngAVtBHh3UvUBNQ7wFuFo1QDsY+0
xzBActdPTE+YJcx/L/HA9adI2cw7hmtwSz2AtHgL2b2V27y/9elvPAWyoeFAshkM
rK43I14cgtgHkjKqSdu25/n2wtHU2pajfW55hiWrKyJ4xUxOINV1cbYSOyj4fNNA
WtrXZyZDhScJz+wXkjs5h+PvRI5UmVFPZz0+3wpdRXJL4c35bHfe8jV7MSZ2q+2Y
ls56pLlP/pvCMFtAtDZOa9g1Fc9mNiWLVsi0YHBteZri4iplDvw6xrYwn7qFXMJ4
XCBg3zpTSi7iyJSvqcrUT3s6fj+MsBUH0nPObmDOa0TYi/OZNI/HYRxWZVpP3nmt
GzBK1/SUbdv33Hd/5GAEb41NK6SFwfZVqCy+vJI8Yt8o7dZouO4zggcIQv4Oco8u
wj2OeHxiGvhImXo1tTM1zidLsdKoLpq7B9TqCUHtczpzCdQsgvSWElzphb0xmy1E
0WTYpXCzNrFiqm/KZF66qdWwx7MPQm5qktMvtUfRm10fvZ6B9uI0n1aGbe+E/YLt
F9peE/EJGQNfrmsPUihE20ibWNWXY/fo7d9kzmYlT/VKYJlcBzkHDnvBCFpM/nLt
pkLiVzZZIjWThK1dYq7yQOtlNDyDT3FZ0y4ixYfnaMiv03H1vXL/nzgzYJdTZV2C
3cOkoAJNO4q7yU7yMS6jB7B3uNkwgtJlUeEPFqIzLbM71AtiybsXiktc3QO+b4dX
TyKiGVVeC4Tuz+g+JfeDnXqw0LJ5sHmrWW83WWckMxS5Ley/qudr8F/l23wcmN8L
4uAb6yHHqVjxmpAFZHS3Y7H3hfPVyM/Is+vYG66izZ0XPZcnFKY+E2aP329OfudZ
EnZRTES8VYBRh9So+WIg3zm0hLEYGlHFGI9vfDyeJ/VYyXLyu8eHxvLUGPTvgPSR
sX77uEF8k7b68PpmQfnSOys389VZQPcST4MgsslQMcOaeQ95Vtvi6Xc/6AdQtvPO
21ZfkaMti3qtVu4K6zNMcgxzBpAzKJ4TdeI+q046h5MvYXx3+jrU0wujixxThVHa
EJ30HrSImhJdL80560/z7RY9YkgoNhcMWTipmZYaZtGE64X4J7QUK1LFskYtBMvd
JSqloL84aMJIAhS0KfSu/K6Ha4XzzZm4kLVDR4T0OTSsxa6iScZF9xdsAfMEfmeU
3P60Oieps/HofyDfIMsPw48kG/nYsMU1nLIZCkqvHKYP4/zrc9FLg2VR+fgng3FL
si803tr8wAZcFdl357PHrJUKCJIylRf8bDzjlkpHrHwq+Qjo+QB4OHM/Hr8poig0
0MBsFfxs+a4CITlXzgViohW+1cgo6wqCwWJruljWox+3+2PtMUjegR1ZIncHUPJN
LmNRWBPTxar2aAofd1pDgvoIlKs1vrk5/5Z8VXBpOYasVNo7TTkkngD3zhoaMdl0
3cG/oj2Mz+iD5ne3bWaUA3zayPZOh53A/JdmdBZxcVO9ojOwGFIwUy5OSgH8BCgV
Kdr5klZfuvgQXlMftKUu1O8cU/eMFEKXWYtuqz/qt2oFgBIHWqA/MfmDH7qMbHJu
LTZfbnaWn83+2KtV5snLN93rZXo5dlBRCRX5F5IncrXjoDlYO+6awPgA1FQQkPnE
4ggXKgi0+NWaAJ6GpGj0u2akyxtooo0iiOLa6qC7PamHuer5HBvqguJLOUrFwOMN
DPcJEE5Rnkj0oiyvFVsxf7sj5qCfydUH4AqrONIy5SDgXiOXmE/9mfIFRJWncNEI
AJBvyU0Mi2ucGaXdPaw3AZITuU2NieVQXPAz+Y7z9B0oo2ChBKVC/Wa238A2Ebhz
2gS+KvAI28ZB3Fjf92pzJL1I3ZryOQFjd5bUqM1j2Xmxr8iRairSlTFMK+0cxeO0
Wzuqj+zL1kwQ0uPByfS/1WcYyxDH6VVx5hGT+pTtf/qaDsa5Gfjr4tt1mG/KSjPc
lVkpEzgdlkc9P2RV+41cnvvOCzf8klvFxTPUH0r6GcZOP8fE/Ml6dr8FNQMrV4cy
OwFZl5SeUrvnkhdq/KPiLVhZ7jfMr6/958DP0t5gNdBhRrngKdyxCk3Y61KrfgB9
y1b7m7KoqHzHXIRwMx9CmXmYQrBxWOaS7jXxfED11gHg4MCgnih2BG7e8V536qJo
sZNJJcndeQvQJJ80JIgByAZ3IZw+S1uzMwG23ROkFIzAeyjsRts70yB8JMVRhbIF
pUzILg1ugxywnakK7bnMLRZIYq8mCE+OwzP9OKELuBQmXc8bfPvIq0i/yoc16aMG
k2rwa8HmOJus9p8CCrsMPjtzBUTDrii7DffXvix6Do5t3UHnNbGy+gN1PUow8qSA
H9LvUl3X2u7hO4lgYoeDRmmZJlqKYx+fxg+SCXiDOSdfhy5I+wPkZtXjBST7IwEz
53QKr+HyO6KND/QvoEIvoZmsBRnTGYzAXY/UAhGdlpbYb8v+XBHw1ZG+soWfbY8n
ik/VtRqb6feVwTawxlWigxWGWDo3ao91evQ17a0q98yA2hU4rZGRC42hXe7iMH94
JfFFwy40b2In9SaKtPO+kxCW2G8Yt3UD++99Culox3W98fXbhMG0N3N1Tc1+5A2r
5C3u46dgpo1QZsuL+ZZ+x2Ft9GLuDutboIn+1H6ASjgcEtYR9olL9aY87OycI8/v
y028b4bS9uuG1aPxODOTXfopslmKWGtTGZyxd/OuB7bPFDfDNzIv5SdcsYnzNtH8
tPUlLUdYbwaVd5cYeF5ZkU7vzOg5sUtnjzdwXclC4pqcbp7WadKbaWzaQdwWGM++
odow/Q1qqG7OXllaJaGnnbVEb/PZeWFdfQapgNEWxCIqR7Egle4Nsgwcm8C6rtkC
Ub1niCh7319RnU0D/0dCmGQEwylS61LPfmz8yIrqUNO9tsmf1EiFBvkkgMQg3vc9
qwWfYcAZaaoT2Rxqc/P9fb44B0mpitLkzswjU+Hykcmcqhrn3krXVE1ASedYopPT
EqfkNujDDrXc78UWDbRWiFO8DE7vBHWpMSlfPWirZXTVedeh2+xIixDfu7Halhsm
6mRflo/MXShcJlYElB/FrmG98jGB2lXq+26Y7llAjWif5yBe4GtRSA/muIgufOQM
Lr7d+/vbRPIsdcJWdbG7eGC4QXUzF+Y1Meq3jG/iwDUOb21H2zjqxsNpt7/rI9T1
SN4p4fSnoFx3EpbN0J5TszlyyP1Wg3r1K0I1LP4C1mql9SI9UN5zVramrG2MSUvv
LRsWBIcdIwDT7wOPTYKwZRAuRacpfYKcqkGQ+UPe13VrAxdNcS7Tl7sVM6KOq4PR
OMhHv+eg0enIAqjKJ8yf4uBzk3y/C6oQ/+dsQFSyRoo0OJj7bEIjD2znnGY/AcjK
+Bq0vUNGjP0iJX2MmJDu+OKncl57RFPYl3Vv5oqGz7FFKndqfgHr/15kSIWy75Sz
7rpKVFGZKjs+mxo8CwmLs9+1g21NDxm2/ZRmS9a+32qBnBZ06WCi8G7wcR7N201f
DOysdnuaXtCzS36ZOyehYFubLsOvdn+1wJ69C/ItdSOjaSgL1J+0ph04IOsAWNrG
iDThqKj1b6aNkxh9hTgeQnEOQeYhVKj2dvSNqh1pQbg6EJxXuMSokN/5RM7bAlCp
rzh26CktDllntxRdZSKZ4VxmOZPSMwM8koHscX+sat+5Vl2IlJGw/RGyiqkeO96i
oOJvTsC3hep+jL2ikHKcpKV5ccfpFN94ONax4VIPX2qImVG/z0egz0qvEVuDmQ0+
apJwy0nV13dHROv/X3MDKbRCZc/848OUGpgIzBmZ69R/f5qyiFfGGKrKl2w9MP+T
4FOL5CVbSkvF6Tw1eET2reJKl5em6Qlv2Ih9TcW0YccQJUfnXuYzwiBMNUetmztA
lLI1qs3/QrSlZPuFI/hFfqFDES5NTDAL5hvyKX9QwNwAnh+Uv6FsE84pTcY2vAhK
WglhxKPtaP5ri1gNlefLLiLe+tjw6aVu+ztoTCB9jTFbyMr2n1pvVa1CmTo6l7lA
mlsAe/nesoxMmn5rQUlEOfSfpan1/7dh89UOTeGB2bZb+EBuZ29v7yhkyYm1oluL
CaoLE2NASMogblBs2XjkAzSzccvUIYLqcKp8QrrJ5NAv+C+VG+EyBHJCP1l6DCRL
Xrf6/HwIXmBCcYDopnOj5aNdaG1ienbibB2RpHGlrY4rfHtFDjI6F2sFIKuXvOgh
fVDrLum1xx8+MjLIp3u+PoL8DICCYHU4yawAwMoXBo6MtBITggySzV/78OjGW2UA
1DzEjQuGwbYi12h0qecQiW6xJTfRnu0u1vFOLT1wP17jfzP6HRPJF4lLiUbkPfMr
AO+XpCCCopCI5VJyLHliBsx27sZg0V+Agze6WFponDyIH3CCH7uapYf7gsV5krbl
ayUqPTPcG9+OhDjZPU6mhGKZGU0Cv0C6MCXivpi6478sMgWNd6nHmiKBK4jW07Kv
Aoq/jHWCEjGpMOFQgx/LIR5FS2lV730qv6zNaKi7inDud2rJBouZiSukkiE9X3y1
RFJvEtcP76TUHDKoP94EawLq2gg2ys8pfy1askrDPForIEmS+0G74ISZc1B150Tn
TCAyMDKlqMBt8xvPhrUfCEd8kwSnpAK6D59UStup8EIgBVwnbM/wWSzMK9HkCfAp
FZe472V+Qka3vZVonSXr1E7vmZWfH6Vzh+KiuFMc0h6/SO4m1nODeZO5ef1KaRHh
2vBfmZlxTGSgdj/R4lBOenkHQGOPaibTEIFbD1cwaBK1oRo1iCcYK+JZcBsHMOip
jtTnrsy3Jgx2AQR4lehJSb7wul/+QoQro4A3EQuLtVIn5uUhj7h8kiY200yZwrUM
JYZ2aX+/GkezgP0Uti3LecpiTV6aZj2Ds4RVn0eqPGypPTEcoM9mqJ5rK2pF+UZz
JkBRte3a/HnB9NfUR3uXIFzIM9acxiT9Nj3WyVkH+lW9Bz2nQvrYxfwv6oY1L6D+
yXtFVp8j97yPN7sOFpjgk1txN+mWFkrwqobqxtvpe371quulkmWkzn0jWlAh/OsJ
XapBZrWkmgD2kNlZamk4gCK0Tq4+1K+rAp+RwVtxDCp7q534SaujI3dIaACGmzlC
+IkPQsS/jyanFHy7xVv4LEfMGXBgWrPk755pbkDNi202ec9GZz7tfYa/loro/2IE
41PzgnUGiuABiiy1dL203W4T4O5c+PQ1zLKOvwgX/x52GP33CwbeUsGwkYteJnxE
Hy94xUEQ+5T4x0tUC25KkIcsSIrvxooJou1lfxJPWkMfo0mBhgMFtyT6k7/lhT1K
zujOh393ciUs+syWj+Z5oyb1OtwQU7xvUvjiqx7pfgfS1geQb7zOGAAJuCWuo/sb
WKrlCY5FoF8yTQgFJAoKuW46xgPvrJnGc5z8I+L8cHAJ9ejP7q2OWpBnBcv2xI8o
PA0cw72hWVYr408aagFnxYUR1L9TCQfK5pmiKtGqSiVHtxPGpa2uHnFW2W6pQB6D
g9gCOsFv33goibEp29t5iPBSQsla1QP4V0FT1hNLqstGT9jn2QlCp8C42HClv3Xd
O+VQvR2eq+OWQuA1BPu8mfMDXpp7qDwzaia7D3H5IEhbPPlSUUU4pOJCU0srMDmg
relb6IMv8HjbdZ3mxSHhOR2yFFVe39a7rDZZrG5/dcrpZXHXeakdwvODE3ONnBqB
0cHc9edzIMYSQsAapD+X3+Fif00YNHH7dK86UFZ/V0+lrdvETDtjgITDqBItOVoZ
/8BsrsaA2Jx8fvG2SHdO75i9UOWqdbb0WWP1ccCr07Ba41ZobYkPL0psed9f+p3a
BdQFvBH4zpGP4Cvy4nDlJUFqVGr/I2zbgUjpjigziB7QhIrwBgcokwHJDunOaPGg
eaqvSd8yuCz/sCoAcKvSz9rG6iQilS+3q4DxBWBpmiE5U3fqqIifHUQEpCV/32k2
TecV2dS8YUgdWv62F5X9aubzOkQBQNftFQPohZdX6o9E6f+4GNf3cdujMKG7d8ja
9TibD1OaQnBtY/7EjVgw8Vei/XUgnHGLIcIQxJITiqguKQ3tllouNpYsHTjuRJ9B
VNDuo1w9WB6NI+JieNfhDwKlIrR/W3lAFWtp8a+YT4V1PVTbJ1Nk3JKAqeispDTM
/q/n8p/jrE8WBtDchEwOvgS5O/oqv/L9kyC6HGE6ki1pr5k+TkttHCceCcUSjytf
Cl0d8mBNxdk63wxzILY8vkYft9BZKkvxxk/ZeYW64KRwA79X9qPOIuNS6yeFZvpj
7WjwoScKlXfNFgANw/jNL3Uw9Q8uzs+3FtNcDk0LdXcVOeTEY1wXI1Fl4KqEiS1J
ohdmVrfeiFWzltLiOckv+Dz9HDe8IDQPdV4JcFmcM3qL0QE7eU3m9zBEzWwrlOBf
8xxR8qrKABWatd++cni/jJUvxHvi92GnTWLHEGh9t42Y4ty2jTdMnJbmTn1IfzX/
b/AgHFYYwbswxlMKTeQttNko9jrL/2CFXwmh40XCVkkHob523/Nj2MWaD+IjY8Aw
Hj9zSgdNovpx8d0EiYJLQdN9kHkShqSpeWgfDgfMto+gUCPK1uwRNBX5az7rhNA5
qmMCJWv2bb/2oi7HW37gkheMOpmKaFkCH//Prt5VQ1dYZ2cj5ZdniVaX1PbfbPxu
MDufn36BrUDlLDFSqL7N1j5cd+82O2I8I/Lc+zh6ty8FWh4LZw9N4ThynUyb27iC
D+8RSVN+rsN1MJALQ8NKJY90wuo3Qip6ubr5ioVfrE4RDs3/nN8jM2tVvnKu/b4x
f04YiZwbRoU88yQlA4ROp8glh7MpA7gUfN+AgjxNhdKOE+ksHzXQK/Q5jEeircdO
jO74ymd8lw9UTnuw5jhj8oJdZ0THRO1o1YbLgNiQ7Z8BINHgEYMK9dv9WtTYt7iZ
yeKIopdCnmnXmhH5WRzr2M7C/AIjz9mLbPgpd3yAdKPziFABHr0Swgkw7JXIWwhV
OKHxwi35Oeu8h/RZcH6lAX9maafIYjk80DBl78pMkoTKtP34PWky1dlNNxaPnRAD
C1iHtxoMTooM/gYhLdec6UDBaPm3vGxE+QPezgRgOvAtwC+9ze4MdOFUGNjvRjAH
ksqqUurLWcX19mVuODw6DxSZ13yuloabaAMHTECal74nRzPYuvbJGhTWRQQ4Ke6Z
20qyUV3L/LOvqLE7NlUBF1WKt8zYm3kA31TqhYa072BeYUNeaJE2Y06AEMYX43gE
z3TinnIVYy/ymtCByAiBv3lyVPAl7G3qhKDTuzaLMdlzxJmG6zvB9gC4nN1VL+S9
6zIxAqWAbE03uAd8zpc3IA4EVFOxyuNiN7G3sLwfE4bf2jGmmmNOg0sokwY9KdTz
B4CAW5QydHyrvs3Bro7hscg18Lin5XtceawZfWfdNybF4zNBShzVnsIpoyrZ45Jb
`pragma protect end_protected
