`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ArynLiqH26XKWrqnGnNodDxZjQZDqd0CMnrtsynIZX4gklcQM51kPExmml+iTLDL
YxqGrHzmaZvMNFwGOmXwnlCkbBT+fpHgaVodF6/DOKNxPTLKR6YQhzg5pHDRq6dK
9qkHOJNTTgs+Cgi38+FxoZWGyd1VhO/O4cG8uFhwoIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
A9PAab/0UbtnwNu7mQsRAGylKZUZZ/6YUa22jPTKqMiC05GkDM4Is1GyeUSxuXv9
HPh0vHQMrtyaqkVdLbVocUDsMHBhTSQyrn+FBl0+VQyzX97IIPy6zT+jjtjaqXH9
nvRMQIZK1bOovabpJkMDcBJQJs6e4tkxLgVcdyoI0+ysL9QKq1VaVCVdXtTycMb+
2zLjw76tnQsUgNWRX4uaqRvDBJh4F6MPazyLfZtH9KJ/1cK/A1uoMNNy2ciugLL2
mWpD9KmJV9DglLSZy5jplqby8+eEp61PQ4jOMjVOM7FWgG5YVnZ03UZ1GXdNmBra
ALBH3jbTKXAIyWzlIX4Ay8hu3aixHUmDfYo+a/xR477Q+SZRNN9ESncfxd1T2pI6
vOJw0YWbhaS85xl5mScz80gij4IszsRg1MNCZWueMQIzXG9A2k29pURhO/GcMzDi
/EnBtY88gDGJFsyj1rD1dLDvjbT/x3cYegC9JZPQr9RZ3rN83QSRX/i8J/A83aXN
ix06uOxYxsorEvGvALWzBYaBKuTtgp77DHZT52LXeaehLr5oGf73Vxv/TLj3X/pX
Bbw2i9570IvAbpbcYRvCntQ3Ef2kfn9oKk/Orl5x6+vmJ+yisWMZ80iaHN/emvvR
bqB0sEMh6sI57Ie1ORxUasHdFVyu5HHa+vTC61/pPsY4UKSoYROHMrdhFRfhlxMr
LZWMiYkM4lKzukYipfItrEP/cUC0rr9cYjGdDSh3wDR87xZo0wdvaZcXUPZKH5u3
ACtzeDwrrLDi3Y1jWIRdKPycxaXq53D83xhaGOZwLAMOnykLE4ffZ7VCF2UEGpDf
0T+SFgQskK/petV4f9LBHNJi7Yxm/4jIzs3jEfo1Fes488CFPN+586MAaJf74PKc
ZSsNiC1JN1GzMBXDGcmHlQKSmS7sJ+hfTHLlpa9stzkL7RcoMKS456xwBcUU9jmh
JyJCupKp8HHBkXbJkIqO+cJ0ybsFHGrOo/ax+layXdEmJ0CKuPsacdKVxaWRu8zh
0yGPkl+Dn38Nqw5wWm0hUJu/ogXs/+VVoyhMeVjM7WD3PAsJ3GJlKds7ZiVw1LP1
AZd1MyJozPOnesK9bXCGeT9wP/fc3Py/PyN6j6jvXKufNA+u32LlcJJiL/v2ylgV
gm4vC+2haBaIy/7XF0w3ihstKDSLGHrtvmfgB6Wv04BJRmNy0ExilsNEraKTRKwr
3565Z2Nr+xuaV6iMOeMzQLPzGQP7L7mq344ZM5X7Y9ay6qNP9z+NBdjPcnRri6HP
vyewmG5N9xdshhP0yiOY5wQXAT0YRF3QOO676BAvEWWM8UINsl8dIk8X7DEwyJvm
JwllEgNdO4AARJbX/Nxwah/W9WoyeFjjKXK6pyiZtwjMMdf3iZRnPkfVZn/+qUYd
jgprVLvT2kSLnLV/K2nU4/l6Obfwv5f08wmFyWbSvhGasZf5gpfy2ZNpEc692+45
mIsJfousZRYA1zMB4l88nDsvG91gj4b9M0cflnkzLUHrcDOqUFInBq1eALB7MYoH
cecFLQItCOiNLTInBCvH+gSrusxqvhnQgsUjB5FUHik1rZt+ykk1DBY4GOhq5qkH
v1ZHUkIoX4USI5hl/XxLvhqIiAUMeImsq6l18acTl4lhb9doiNtEMAXpO5aHJYGB
tg41W7SuxR5i0WNfGBe6SjxPc9V1vk9sbLaez5DIIOEeVxj7IYhVtHMFPc+gDLKr
FITaGtFyIa2/tKv1nGS+vW4o8jHGbGohpNrIXMp61T9iwJr0Mn0Ds1wBh67MgIz9
izgwBwcwVzKAGe+SuZ5z204kOTlaO60p9dm2IQXUNi/UIbcRuh0XcRbVIRUENlxR
6S3V0Tw+Izu1lcWCUf+XNpOOj1Czehnepx/+PuhSljXqgCsyYlrUAiXxzUGmRzBz
NXXusHfQ7DyV774qSqefTHH9Zp1u1yH6iNphzOJQMZ3OxRDmFS/CAVouhWcNhe9g
TMFB2UjJ4JqkzI8APZyKb3aMHCn5ISzjSgXfKoum6T5PNqHPmT677kgsQIdzni9J
ur9jeRwq9jHGerWQLo+idJycOcdXAmfCfnkr/1GACoyjR/i1Ns4lXWjioj9eL/af
D+1iejrvaae05Fx8+4WMvbmG9+0ND8v6ySyecEXbffsYVPTyZpMUwiJeRQxpztD+
yykQkRjZuvivAgCVxamuo//rcZpOJseM3H/s88W0CzQ4U6ZLRlj1oM7slLrT0iD7
pS159sFcXX4NiQV/k4q6sqOllmILSnToe6UeqRNLwBUElp95Zxdi6Gk5MF31xFoX
atqqjwwVoGOH7kg5Yk4o1ZFCUQfo6fq62gd1l3nbZNBgI58+sQybLMAXiskR5taa
4++MuUAF2Fdq5zbQ0MEJVisW504tj7i+AswI+hEJwzvD0eL6RrF3vULE7qphdKlh
nS/fhpeJst1YqUSbzpuX0WII3S4LQQ3mgJwnUskSAVHEHPVetMA7reCGToBr7/d9
vLL734ki3MweJPMxf+T8MyNa/oBByB0yZYZX8jNU8K5IMWBYtVXFs8XTmkBDvYh7
QfLX7WyKmLqwa2vveoBbe8MTXWkby2YW4ABXwd78S5RJZtU49G/nES3muw3AkU3q
hz44Pmt4SCvOmvMB9qG1HdXRla9AhNsDHHFiA7cFjlCYr5OH41W8vfAJttdTCjNt
8q1zj+ub4qxZtREEY/1xe/y8DAOovZU6eq4AY2rFrJbvdTXSNllQVNHh5W2uLOUS
YqCus8pOwJSz/PGlbYbmiMVYBl94rTYzwmUc5Ee00c4U0RYXStCDEVCavJHfLG++
yJcvEoAL1pwFGby5HrTa5HBVS0+aedXWG76w/oSrC7zHi2mInGiJPgcOJDEiQj6r
gijnFHfd7g0lHkPRc2iuWJgDqDRK2XjMFXa2hwQcAZvNkSaqkOPqxYmpExY+CaPR
KwZeELzLIvdqp0wk6JOYN17/mFcm+NBgMn1ij40MLk5uV9vaa5NkmcG9JV1WxSnQ
/45JCbC9WZ2pYEg0vnIT1W8wdLTn+ZcC4qE13R5CP7ocPlRY3Wqw8pClWDAbsnbl
UDS5whIqNHFQk4Q3d2gArg+5K7jMn4/t4Kj92qEcyKmvH0vsrIjgFtMZMoVs9NFs
+wIEBVL9U2YgfNeooywnX/+SOA7mpAsL3ccYDasId1MiUKEOdbvBXRHv13u+vjU2
f7OL2bSZoZeVjSUOok4fVL0Zx2vmH6rIBR4hP3h1McWIkBV8/7zGo/9dw0g8XM1A
ceqUOJkhHfArkNhp7HD99kuiecmWQwnnAo+yHVagdtKS34gKtb1cM1EIZNGACHD2
k4dnKkoTe41BUxJtiZ07/RU5jQ3RLYEMsrfxRw+L2hmZKvKG0ckFWRjwm8ZKaWA3
upbnXbSiI4BxKO9vFXXn04n8Z9gOSuRhY2XcQ2wdlfUixN1tJIqK8stcamNCRKTz
mCFmOpjy2b/9H0Zd3RfDKxIIpIpxTQuvnvwZad9IIk25oHngPy/lt0+PPlrdfPxC
M5XwSvvxtGVNacUIkXR4QDsGvMJHQkdGUUYGIryRrCpfymRHdKbhtViE0sWHCZuc
GnaxJqve22+NdVfLnkmNzTzi3ihW6C0ORVfFz+tH5McjsSUcupJwIoG6ADuwPXLg
hG1nSjJ4uPNQ2JW8YsL1nWko3KEHxGgJ6RvrW9fCiOz4ZpYrKU4W2kjEBa3cz6Tt
t/xKZsB3W2uxc5t2M4leX2VgZSFUV1fSS4Oe8kvMsetLCnm72BfnaM5fqQBELyE7
2JTdL8pX6XQCxreGcpRkXbEH7vJxv7Ty/4HJud6bEyDhLWOqZcMrFT+LMTYWtzSl
YWDjSSaRM9meElRy4KLa2i2BFeuBcsr7R1ZNCc+Ap1RprNndNL9tB1chAuqGDCrt
KfI9QFW8F+6n0rJVEy/imcsobvx5BlWMNfy5xsk1di3jDfvVp1DvVpttk2cmYUqn
+eYjVZubRCNz0EpzHi2i61u4NBKULYg1ekOXSOthAvh0DLz9idrFTHfPcjG+wS2x
p5E4YFrRdYRRzKBkJGHbBbfBWOqptGJnBYBT+V1RIZ4+EmWItrM6r+u/wRVIHdC3
G1hl2OuCTc1OmhQN5xvsKcsPTNal2lnau12GCaLanhRrhBG/oeCFKV7W1U+T9AxZ
jY1BxBr2qxkv3htj//RDHA8TQ9Tyc3E8P9+xsXLXi3s=
`pragma protect end_protected
